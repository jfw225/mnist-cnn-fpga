// synthesis VERILOG_INPUT_VERSION SYSTEMVERILOG_2005
`ifndef __LAYER4_SV__
`define __LAYER4_SV__



`define maxpool_weights_JWCVA parameter bit [15:0] maxpool_weights_JWCVA [2879:0] = '{ \
	16'b000000_0000100110, \
	16'b000000_0001001110, \
	16'b111111_1110111010, \
	16'b111111_1110101011, \
	16'b000000_0000110000, \
	16'b111111_1111011110, \
	16'b000000_0000100100, \
	16'b000000_0001011111, \
	16'b111111_1110110001, \
	16'b000000_0001100011, \
	16'b111111_1111001001, \
	16'b111111_1111101010, \
	16'b000000_0000111000, \
	16'b000000_0001001101, \
	16'b000000_0001000000, \
	16'b000000_0001000011, \
	16'b111111_1110011010, \
	16'b000000_0011110000, \
	16'b111111_1111010110, \
	16'b000000_0100001000, \
	16'b000000_0011111100, \
	16'b111111_1101010100, \
	16'b000000_0001000010, \
	16'b000000_0110100111, \
	16'b111111_1111110011, \
	16'b111111_1111001110, \
	16'b111111_1011000100, \
	16'b000000_0001111001, \
	16'b000000_0000010110, \
	16'b111111_1110001100, \
	16'b111111_1110100011, \
	16'b000000_0000001001, \
	16'b000000_0000000011, \
	16'b111111_1101100110, \
	16'b111111_1000111000, \
	16'b111111_1110010001, \
	16'b111111_1101101111, \
	16'b111111_1101111111, \
	16'b111111_1100101011, \
	16'b111111_1110111000, \
	16'b111111_1111001000, \
	16'b111111_1111010011, \
	16'b111111_1101101000, \
	16'b111111_1111100100, \
	16'b111111_1111111010, \
	16'b111111_1111110110, \
	16'b111111_1110101111, \
	16'b111111_1111010000, \
	16'b111111_1111101001, \
	16'b111111_1110011011, \
	16'b111111_1110110000, \
	16'b111111_1110000110, \
	16'b111111_1110101101, \
	16'b111111_1110111000, \
	16'b111111_1110101110, \
	16'b000000_0010011011, \
	16'b111111_1111110111, \
	16'b000000_0001110101, \
	16'b111111_1011011101, \
	16'b111111_1110111101, \
	16'b000000_0010010100, \
	16'b111111_1001110001, \
	16'b000000_0001001011, \
	16'b000000_0001000111, \
	16'b000000_0000001010, \
	16'b111111_1110001010, \
	16'b111111_1100110010, \
	16'b000000_0000101011, \
	16'b000000_0010101011, \
	16'b111111_1011000010, \
	16'b000000_0001000111, \
	16'b000000_0000100110, \
	16'b111111_1111001010, \
	16'b111111_1011010101, \
	16'b111111_1111101010, \
	16'b000000_0001111101, \
	16'b111111_1111010010, \
	16'b111111_1100011111, \
	16'b111111_1111101111, \
	16'b111111_1010011101, \
	16'b000000_0000000000, \
	16'b111111_1010001101, \
	16'b000000_0000010011, \
	16'b000000_0010000000, \
	16'b111111_1111110100, \
	16'b111111_1111000001, \
	16'b111111_1101011010, \
	16'b111111_1111001011, \
	16'b111111_1111110111, \
	16'b111111_1101101100, \
	16'b111111_1111101011, \
	16'b000000_0001111110, \
	16'b111111_1110000100, \
	16'b000000_0001000011, \
	16'b111111_1101111110, \
	16'b111111_1101111000, \
	16'b111111_1111010100, \
	16'b111111_1111100011, \
	16'b000000_0000010111, \
	16'b111111_1110001110, \
	16'b111111_1110111010, \
	16'b111111_1111111000, \
	16'b111111_1111001111, \
	16'b111111_1110101100, \
	16'b111111_1111100000, \
	16'b111111_1110111111, \
	16'b111111_0110011010, \
	16'b000000_0000000000, \
	16'b111111_1101111010, \
	16'b111111_0111011111, \
	16'b111111_1111100111, \
	16'b111111_1111100010, \
	16'b111111_1110101101, \
	16'b111111_1111010111, \
	16'b000000_0000010111, \
	16'b000000_0010000111, \
	16'b000000_0000100010, \
	16'b111111_1100100001, \
	16'b000000_0000111101, \
	16'b111111_1111110101, \
	16'b000000_0000010101, \
	16'b111111_1111110100, \
	16'b000000_0001010011, \
	16'b000000_0000100010, \
	16'b000000_0011011010, \
	16'b000000_0000101111, \
	16'b000000_0000111001, \
	16'b000000_0010011100, \
	16'b111111_1110011100, \
	16'b000000_0000111000, \
	16'b000000_0001100001, \
	16'b111111_1111101001, \
	16'b000000_0010000011, \
	16'b111111_1101000111, \
	16'b000000_0011001010, \
	16'b000000_0010010010, \
	16'b111111_1111111010, \
	16'b000000_0010100100, \
	16'b000000_0001011100, \
	16'b111111_1111011100, \
	16'b000000_0001010100, \
	16'b000000_0000010001, \
	16'b000000_0100001101, \
	16'b111111_1111011011, \
	16'b111111_1111010100, \
	16'b111111_1101010110, \
	16'b111111_1101101000, \
	16'b000000_0000100011, \
	16'b000000_0000001101, \
	16'b111111_1101001100, \
	16'b000000_0000110001, \
	16'b111111_1110011001, \
	16'b111111_1111100111, \
	16'b111111_1110111111, \
	16'b111111_1000000011, \
	16'b111111_1101000101, \
	16'b000000_0000001111, \
	16'b111111_0111001000, \
	16'b000000_0001000101, \
	16'b111111_1111101111, \
	16'b111111_1011111100, \
	16'b000000_0001101001, \
	16'b111111_1110111111, \
	16'b111111_1111111011, \
	16'b000000_0000111101, \
	16'b111111_1110101111, \
	16'b000000_0001101110, \
	16'b000000_0001011110, \
	16'b111111_1100110001, \
	16'b000000_0001000110, \
	16'b000000_0010111010, \
	16'b111111_1111011011, \
	16'b000000_0001111101, \
	16'b000000_0001110011, \
	16'b000000_0010011000, \
	16'b000000_0011011111, \
	16'b111111_1110110111, \
	16'b000000_0011010111, \
	16'b000000_0011110101, \
	16'b000000_0000001010, \
	16'b000000_0100101101, \
	16'b000000_0001011011, \
	16'b000000_0100000101, \
	16'b000000_0100111111, \
	16'b111111_1111000001, \
	16'b000000_0101100010, \
	16'b000000_0101001111, \
	16'b111111_1111011011, \
	16'b000000_0000011010, \
	16'b000000_0010000111, \
	16'b000000_0101101101, \
	16'b000000_0100001100, \
	16'b000000_0000000011, \
	16'b000000_0001010101, \
	16'b000000_0001010011, \
	16'b000000_0001101110, \
	16'b000000_0000110100, \
	16'b000000_0010110010, \
	16'b000000_0001111001, \
	16'b000000_0010001101, \
	16'b111111_1111010000, \
	16'b000000_0010110001, \
	16'b000000_0000111001, \
	16'b111111_1110011000, \
	16'b111111_1110001010, \
	16'b000000_0000111010, \
	16'b000000_0100110101, \
	16'b000000_0001011111, \
	16'b111111_1101100100, \
	16'b000000_0000100010, \
	16'b000000_0001101000, \
	16'b000000_0000100011, \
	16'b111111_1111000010, \
	16'b000000_0000011001, \
	16'b000000_0010001000, \
	16'b000000_0000000100, \
	16'b000000_0000010000, \
	16'b000000_0000011111, \
	16'b000000_0010101010, \
	16'b111111_1111110010, \
	16'b111111_1111011000, \
	16'b000000_0001001011, \
	16'b000000_0000010011, \
	16'b000000_0010001011, \
	16'b000000_0000001101, \
	16'b000000_0011000101, \
	16'b000000_0000010000, \
	16'b111111_1110010111, \
	16'b111111_1110001000, \
	16'b000000_0001010111, \
	16'b000000_0010010011, \
	16'b000000_0010110010, \
	16'b111111_1111111111, \
	16'b000000_0111001000, \
	16'b000000_0000000000, \
	16'b111111_1110111101, \
	16'b111111_1111001111, \
	16'b000000_0001010010, \
	16'b000000_0100010100, \
	16'b000000_0011101010, \
	16'b111111_1110110111, \
	16'b111111_1110011100, \
	16'b000000_0001001111, \
	16'b111111_1110010010, \
	16'b000000_0001111000, \
	16'b000000_0001000010, \
	16'b000000_0000001110, \
	16'b000000_0001011010, \
	16'b111111_1111101001, \
	16'b000000_0001011011, \
	16'b000000_0000011001, \
	16'b111111_1110110111, \
	16'b111111_1110000010, \
	16'b000000_0010101010, \
	16'b000000_0000100110, \
	16'b000000_0011000111, \
	16'b111111_1111100011, \
	16'b000000_0000010110, \
	16'b000000_0000010111, \
	16'b111111_1110101110, \
	16'b000000_0001000000, \
	16'b111111_1111011110, \
	16'b000000_0010101011, \
	16'b111111_1111011100, \
	16'b111111_1110101101, \
	16'b000000_0001000011, \
	16'b000000_0011101100, \
	16'b111111_1110100010, \
	16'b000000_0001001001, \
	16'b000000_0000001010, \
	16'b111111_1110011110, \
	16'b111111_1111110000, \
	16'b000000_0000011001, \
	16'b000000_0000110111, \
	16'b000000_0000101110, \
	16'b111111_1111011010, \
	16'b111111_1110011001, \
	16'b000000_0000000011, \
	16'b000000_0011011111, \
	16'b000000_0000101011, \
	16'b000000_0000101111, \
	16'b000000_0011010100, \
	16'b111111_1111101001, \
	16'b000000_0001001001, \
	16'b111111_1111100111, \
	16'b111111_1111111011, \
	16'b111111_1111111001, \
	16'b000000_0001000010, \
	16'b111111_1111010001, \
	16'b111111_1110111011, \
	16'b000000_0000100111, \
	16'b000000_0000001011, \
	16'b000000_0000101000, \
	16'b111111_1111100010, \
	16'b111111_1110100011, \
	16'b111111_1111010010, \
	16'b111111_1101111011, \
	16'b000000_0010000110, \
	16'b000000_0001101011, \
	16'b111111_1110110011, \
	16'b111111_1110111110, \
	16'b000000_0001000001, \
	16'b000000_0001010101, \
	16'b111111_1111111100, \
	16'b111111_1110110000, \
	16'b000000_0001010011, \
	16'b000000_0001000100, \
	16'b111111_1111001000, \
	16'b111111_1111000001, \
	16'b000000_0010110110, \
	16'b000000_0001000100, \
	16'b111111_1111011001, \
	16'b111111_1100110001, \
	16'b000000_0010001010, \
	16'b000000_0001010000, \
	16'b111111_1101101100, \
	16'b000000_0010011001, \
	16'b111111_1111111110, \
	16'b000000_0011011001, \
	16'b000000_0000000110, \
	16'b111111_1110011010, \
	16'b000000_0000111000, \
	16'b111111_1111111011, \
	16'b111111_1111110111, \
	16'b111111_1111001001, \
	16'b111111_1111011101, \
	16'b000000_0001101001, \
	16'b111111_1110111110, \
	16'b111111_1110011010, \
	16'b111111_1111111100, \
	16'b111111_1111001111, \
	16'b000000_0000100001, \
	16'b111111_1111110011, \
	16'b111111_1110000111, \
	16'b000000_0000011011, \
	16'b000000_0000101011, \
	16'b111111_1110000110, \
	16'b111111_1111110101, \
	16'b111111_1110011001, \
	16'b111111_1101110111, \
	16'b111111_1111110100, \
	16'b111111_1111110110, \
	16'b111111_1111011110, \
	16'b000000_0000110001, \
	16'b111111_1101010000, \
	16'b000000_0011000100, \
	16'b000000_0000110001, \
	16'b111111_1111011010, \
	16'b111111_1100100001, \
	16'b000000_0011001110, \
	16'b000000_0010011101, \
	16'b000000_0000100010, \
	16'b111111_1010001100, \
	16'b000000_0000011101, \
	16'b000000_0001001010, \
	16'b111111_1100011110, \
	16'b111111_1011110101, \
	16'b000000_0010111000, \
	16'b000000_0010111010, \
	16'b000000_0000100100, \
	16'b111111_1000101110, \
	16'b000000_0010101011, \
	16'b000000_0000001011, \
	16'b111111_1100111000, \
	16'b000000_0010000100, \
	16'b000000_0001000101, \
	16'b000000_0011001011, \
	16'b000000_0011010000, \
	16'b111111_1101010111, \
	16'b000000_0010011110, \
	16'b111111_1110111110, \
	16'b111111_1101000001, \
	16'b111111_1111010111, \
	16'b111111_1001100010, \
	16'b000000_0100001110, \
	16'b000000_0001010001, \
	16'b111111_1110011100, \
	16'b000000_0000001111, \
	16'b000000_0000110110, \
	16'b111111_1110011010, \
	16'b000000_0000001100, \
	16'b111111_1110110001, \
	16'b000000_0010111111, \
	16'b000000_0000101001, \
	16'b111111_1110100000, \
	16'b000000_0000011110, \
	16'b000000_0001000010, \
	16'b111111_1111001001, \
	16'b111111_1101111110, \
	16'b000000_0010001001, \
	16'b111111_1111010001, \
	16'b000000_0001110010, \
	16'b111111_1111000011, \
	16'b000000_0000011001, \
	16'b000000_0000101000, \
	16'b111111_1111010100, \
	16'b111111_1110010100, \
	16'b000000_0011100101, \
	16'b000000_0000111000, \
	16'b111111_1111110110, \
	16'b111111_0111101011, \
	16'b000000_0000011110, \
	16'b000000_0000100011, \
	16'b111111_1110100111, \
	16'b111111_1100101000, \
	16'b000000_0000011010, \
	16'b000000_0000110110, \
	16'b000000_0001110000, \
	16'b111111_1001110101, \
	16'b000000_0010111000, \
	16'b111111_1111111101, \
	16'b111111_1101100111, \
	16'b111111_1110100000, \
	16'b111111_1101000111, \
	16'b000000_0100010001, \
	16'b000000_0010100100, \
	16'b111111_1111001010, \
	16'b000000_0000101100, \
	16'b000000_0000011111, \
	16'b111111_1100111111, \
	16'b111111_1111010100, \
	16'b000000_0001000011, \
	16'b000000_0001101111, \
	16'b000000_0001001111, \
	16'b111111_1111001001, \
	16'b000000_0000111111, \
	16'b111111_1110100100, \
	16'b111111_1110001001, \
	16'b000000_0000010111, \
	16'b000000_0000101000, \
	16'b000000_0010000010, \
	16'b111111_1111101111, \
	16'b111111_1110011101, \
	16'b111111_1100010100, \
	16'b000000_0001010001, \
	16'b111111_1111001011, \
	16'b111111_1101100111, \
	16'b111111_1110100000, \
	16'b111111_1110111000, \
	16'b111111_1110000010, \
	16'b111111_1111001100, \
	16'b000000_0000111010, \
	16'b000000_0011100101, \
	16'b111111_1110111101, \
	16'b111111_1111101101, \
	16'b000000_0010000011, \
	16'b111111_1111110110, \
	16'b000000_0001100011, \
	16'b111111_0110000101, \
	16'b000000_0010110001, \
	16'b111111_1111111101, \
	16'b111111_1110100001, \
	16'b111111_0110010011, \
	16'b111111_1110100110, \
	16'b000000_0010001010, \
	16'b000000_0001111011, \
	16'b111111_0111101001, \
	16'b000000_0001100100, \
	16'b111111_1111101011, \
	16'b111111_1001001000, \
	16'b111111_1111100011, \
	16'b000000_0000001101, \
	16'b000000_0011001100, \
	16'b000000_0001100101, \
	16'b111111_1110100100, \
	16'b000000_0010011010, \
	16'b000000_0001001000, \
	16'b111111_1110101111, \
	16'b000000_0100100100, \
	16'b111111_1111011000, \
	16'b000000_0010111100, \
	16'b000000_0001011001, \
	16'b111111_1110101000, \
	16'b111111_1110101111, \
	16'b000000_0001110000, \
	16'b111111_1111110000, \
	16'b111111_1111110100, \
	16'b000000_0001100110, \
	16'b000000_0001011000, \
	16'b000000_0000011001, \
	16'b111111_1110110011, \
	16'b111111_1100101000, \
	16'b000000_0000111011, \
	16'b111111_1111111011, \
	16'b000000_0001001011, \
	16'b111111_1111010010, \
	16'b111111_1110011101, \
	16'b111111_1111111111, \
	16'b111111_1110010011, \
	16'b000000_0100001010, \
	16'b111111_1111111011, \
	16'b111111_1111111001, \
	16'b111111_1101000110, \
	16'b000000_0001011001, \
	16'b000000_0010010000, \
	16'b000000_0010100010, \
	16'b111111_1001000000, \
	16'b000000_0001110001, \
	16'b000000_0000000111, \
	16'b000000_0000101011, \
	16'b111111_1011011010, \
	16'b000000_0000111110, \
	16'b000000_0011100010, \
	16'b000000_0000111010, \
	16'b111111_1110011111, \
	16'b000000_0001000001, \
	16'b000000_0000011001, \
	16'b111111_1101011011, \
	16'b111111_1111000110, \
	16'b000000_0000010001, \
	16'b000000_0001110111, \
	16'b000000_0001011110, \
	16'b111111_1111010011, \
	16'b000000_0010011001, \
	16'b111111_1110001110, \
	16'b111111_1110100001, \
	16'b000000_0000010110, \
	16'b000000_0000100100, \
	16'b000000_0011010010, \
	16'b000000_0010010101, \
	16'b111111_1110101111, \
	16'b000000_0001001101, \
	16'b000000_0000101110, \
	16'b000000_0000110001, \
	16'b000000_0000001010, \
	16'b111111_1110101111, \
	16'b000000_0000000001, \
	16'b111111_1111101110, \
	16'b111111_1110010110, \
	16'b111111_1111111111, \
	16'b000000_0010000111, \
	16'b000000_0000111001, \
	16'b111111_1101111101, \
	16'b111111_1110011011, \
	16'b000000_0010001111, \
	16'b111111_1111100010, \
	16'b111111_1110110111, \
	16'b000000_0001010101, \
	16'b111111_1101001111, \
	16'b000000_0000110010, \
	16'b000000_0000100000, \
	16'b000000_0010001000, \
	16'b000000_0000010101, \
	16'b000000_0001100000, \
	16'b111111_1110010100, \
	16'b000000_0001001000, \
	16'b111111_1111110000, \
	16'b111111_1111100111, \
	16'b111111_1110101010, \
	16'b111111_1111101000, \
	16'b000000_0100011101, \
	16'b000000_0000110000, \
	16'b111111_1110011101, \
	16'b000000_0010010011, \
	16'b000000_0001101111, \
	16'b111111_1101010010, \
	16'b111111_1101110100, \
	16'b000000_0000000111, \
	16'b000000_0000101101, \
	16'b000000_0000101100, \
	16'b111111_1111101001, \
	16'b000000_0001011001, \
	16'b000000_0000000001, \
	16'b111111_1110100010, \
	16'b111111_1110010010, \
	16'b000000_0000010111, \
	16'b000000_0001110110, \
	16'b111111_1110010001, \
	16'b111111_1111011000, \
	16'b000000_0000010101, \
	16'b111111_1110110001, \
	16'b000000_0000110111, \
	16'b000000_0001000000, \
	16'b000000_0001001001, \
	16'b111111_1101111100, \
	16'b111111_1111111011, \
	16'b000000_0010001101, \
	16'b111111_1111010010, \
	16'b111111_1111101001, \
	16'b000000_0000101110, \
	16'b111111_1110111001, \
	16'b000000_0000010100, \
	16'b111111_1100110011, \
	16'b111111_1111110011, \
	16'b111111_1111011111, \
	16'b000000_0010010010, \
	16'b111111_1101010010, \
	16'b000000_0001000000, \
	16'b111111_1111000101, \
	16'b111111_1101101110, \
	16'b111111_1111010000, \
	16'b000000_0001110001, \
	16'b000000_0010010101, \
	16'b000000_0001000111, \
	16'b111111_1110101000, \
	16'b111111_1111110001, \
	16'b000000_0010011001, \
	16'b111111_1011111011, \
	16'b111111_1110000110, \
	16'b000000_0001101010, \
	16'b000000_0010011100, \
	16'b111111_1110100001, \
	16'b111111_1111100010, \
	16'b000000_0010011000, \
	16'b000000_0000001001, \
	16'b111111_1110001001, \
	16'b111111_1101101100, \
	16'b000000_0001000100, \
	16'b000000_0001000101, \
	16'b000000_0000110100, \
	16'b111111_1111001001, \
	16'b000000_0000011111, \
	16'b111111_1111110110, \
	16'b111111_1110000011, \
	16'b000000_0000010110, \
	16'b111111_1111000100, \
	16'b000000_0000000010, \
	16'b111111_1110001010, \
	16'b111111_1111000011, \
	16'b000000_0001100001, \
	16'b000000_0001111001, \
	16'b111111_1111101110, \
	16'b000000_0000111000, \
	16'b000000_0001110010, \
	16'b000000_0001111010, \
	16'b111111_1101111101, \
	16'b111111_1110011101, \
	16'b000000_0001000100, \
	16'b000000_0001000010, \
	16'b111111_1110110010, \
	16'b111111_1111000100, \
	16'b111111_1101100011, \
	16'b111111_1111101111, \
	16'b000000_0000000000, \
	16'b111111_1100000101, \
	16'b000000_0000111010, \
	16'b000000_0000011101, \
	16'b111111_1100001001, \
	16'b111111_1111000001, \
	16'b111111_1111101000, \
	16'b000000_0100110100, \
	16'b111111_1110001101, \
	16'b111111_1101110110, \
	16'b000000_0000101111, \
	16'b111111_1111100001, \
	16'b111111_1000100000, \
	16'b111111_1110001000, \
	16'b000000_0000101111, \
	16'b000000_0001010010, \
	16'b000000_0001000100, \
	16'b111111_1011110011, \
	16'b000000_0000000100, \
	16'b111111_1110100000, \
	16'b111111_1010110011, \
	16'b111111_1110010101, \
	16'b000000_0011000100, \
	16'b000000_0010111001, \
	16'b111111_1101110111, \
	16'b111111_1010111101, \
	16'b000000_0010000110, \
	16'b000000_0000001001, \
	16'b000000_0000101000, \
	16'b111111_1101101110, \
	16'b111111_1101011011, \
	16'b000000_0001000000, \
	16'b000000_0000111010, \
	16'b000000_0000101000, \
	16'b000000_0000110110, \
	16'b111111_1110110001, \
	16'b111111_1110110011, \
	16'b111111_1111011010, \
	16'b111111_1101111011, \
	16'b000000_0000011110, \
	16'b111111_1100001111, \
	16'b111111_1110110010, \
	16'b000000_0010010001, \
	16'b000000_0000001001, \
	16'b000000_0000001000, \
	16'b000000_0000000000, \
	16'b111111_1111100011, \
	16'b000000_0001011001, \
	16'b111111_1111101100, \
	16'b000000_0000111011, \
	16'b000000_0000000001, \
	16'b000000_0000101100, \
	16'b111111_1010001000, \
	16'b000000_0000001000, \
	16'b111111_1111011101, \
	16'b000000_0011000111, \
	16'b000000_0000000111, \
	16'b000000_0000010110, \
	16'b000000_0001100010, \
	16'b111111_1111100010, \
	16'b111111_1001110011, \
	16'b111111_1101111110, \
	16'b000000_0001000010, \
	16'b000000_0100000111, \
	16'b111111_1101111011, \
	16'b111111_1100101011, \
	16'b111111_1111110101, \
	16'b111111_1100010101, \
	16'b111111_1101000010, \
	16'b111111_1101100100, \
	16'b111111_1110010011, \
	16'b000000_0010001001, \
	16'b111111_1010100100, \
	16'b111111_1111011100, \
	16'b000000_0000100100, \
	16'b111111_1110110000, \
	16'b111111_1101110110, \
	16'b111111_1010010010, \
	16'b111111_1110111001, \
	16'b000000_0000101001, \
	16'b111111_1101100110, \
	16'b111111_1101101111, \
	16'b111111_1110101001, \
	16'b111111_1101111000, \
	16'b000000_0001010110, \
	16'b111111_1101010110, \
	16'b000000_0001010100, \
	16'b000000_0000100011, \
	16'b111111_1111110001, \
	16'b000000_0010100011, \
	16'b000000_0001101010, \
	16'b111111_1110011111, \
	16'b111111_1100100110, \
	16'b000000_0011000000, \
	16'b000000_0001010010, \
	16'b000000_0001010000, \
	16'b000000_0001110111, \
	16'b000000_0100001001, \
	16'b000000_0001001101, \
	16'b000000_0000100111, \
	16'b000000_0100010100, \
	16'b000000_0010001100, \
	16'b000000_0000100011, \
	16'b000000_0010110011, \
	16'b000000_0000010011, \
	16'b000000_0001101010, \
	16'b111111_1111100011, \
	16'b111111_1111011000, \
	16'b111111_1111101010, \
	16'b000000_0000101100, \
	16'b111111_1110011101, \
	16'b000000_0011111000, \
	16'b111111_1011110101, \
	16'b000000_0010111100, \
	16'b000000_0001010111, \
	16'b111111_1110110101, \
	16'b000000_0010110100, \
	16'b111111_1100001100, \
	16'b111111_1000010010, \
	16'b000000_0100011000, \
	16'b111111_1101011000, \
	16'b000000_0101000101, \
	16'b000000_0001100101, \
	16'b000000_0010010000, \
	16'b000000_0110011110, \
	16'b111111_1111110100, \
	16'b111111_1100110000, \
	16'b000000_0000100101, \
	16'b111111_1100100101, \
	16'b000000_0000011111, \
	16'b000000_0001000011, \
	16'b000000_0000010011, \
	16'b000000_0000010100, \
	16'b111111_1101011101, \
	16'b111111_1110111000, \
	16'b000000_0000101110, \
	16'b000000_0011011000, \
	16'b111111_1111111011, \
	16'b000000_0010011000, \
	16'b000000_0001000011, \
	16'b000000_0001011000, \
	16'b000000_0011010000, \
	16'b000000_0011111100, \
	16'b000000_0001111101, \
	16'b000000_0010010100, \
	16'b000000_0100000110, \
	16'b000000_0000011111, \
	16'b000000_0000000111, \
	16'b000000_0001100000, \
	16'b000000_0001101100, \
	16'b000000_0000001110, \
	16'b000000_0000110010, \
	16'b111111_1111010101, \
	16'b000000_0000010111, \
	16'b111111_1101011011, \
	16'b000000_0000010100, \
	16'b000000_0001001001, \
	16'b111111_1110110000, \
	16'b111111_1010001101, \
	16'b111111_1111011000, \
	16'b111111_1110100011, \
	16'b000000_0011001010, \
	16'b111111_1110000010, \
	16'b000000_0011000100, \
	16'b000000_0001111101, \
	16'b111111_1100111011, \
	16'b111111_1000100010, \
	16'b000000_0001000010, \
	16'b000000_0010010010, \
	16'b000000_1001000000, \
	16'b000000_0001000001, \
	16'b000000_0100000111, \
	16'b000000_0110100001, \
	16'b000000_0001110101, \
	16'b111111_1110101010, \
	16'b000000_0001011100, \
	16'b111111_1111101001, \
	16'b000000_0001011110, \
	16'b000000_0001011100, \
	16'b000000_0000101101, \
	16'b000000_0000010100, \
	16'b111111_1110111010, \
	16'b000000_0000110101, \
	16'b000000_0000000111, \
	16'b000000_0010001001, \
	16'b111111_1111000001, \
	16'b000000_0010100110, \
	16'b111111_1110101001, \
	16'b000000_0011010111, \
	16'b000000_0000011000, \
	16'b000000_0001010000, \
	16'b000000_0001001011, \
	16'b000000_0000000011, \
	16'b111111_1111101001, \
	16'b111111_1110110010, \
	16'b111111_1111011000, \
	16'b000000_0001100011, \
	16'b000000_0000111000, \
	16'b000000_0000000001, \
	16'b000000_0001010001, \
	16'b111111_1101000111, \
	16'b111111_1101111001, \
	16'b111111_1101111111, \
	16'b000000_0001010100, \
	16'b111111_1110101111, \
	16'b111111_1100011000, \
	16'b111111_1001100111, \
	16'b000000_0000001110, \
	16'b111111_1110001111, \
	16'b000000_0000110100, \
	16'b111111_1111010101, \
	16'b000000_0001111111, \
	16'b000000_0000011110, \
	16'b111111_1010100111, \
	16'b111111_1100000011, \
	16'b000000_0001010111, \
	16'b000000_0010101010, \
	16'b000000_0010000101, \
	16'b000000_0000011100, \
	16'b000000_0001011011, \
	16'b000000_0100000110, \
	16'b111111_1111111000, \
	16'b000000_0000110111, \
	16'b000000_0001110010, \
	16'b111111_1111011101, \
	16'b000000_0001100010, \
	16'b111111_1110111010, \
	16'b000000_0010010111, \
	16'b000000_0001011110, \
	16'b000000_0001110000, \
	16'b000000_0000010100, \
	16'b000000_0000010011, \
	16'b111111_1111110010, \
	16'b000000_0010111101, \
	16'b000000_0000010011, \
	16'b000000_0001111101, \
	16'b111111_1101111110, \
	16'b000000_0000000101, \
	16'b111111_1110110010, \
	16'b111111_1110111111, \
	16'b000000_0000101011, \
	16'b000000_0000001111, \
	16'b000000_0000100111, \
	16'b111111_1111000000, \
	16'b111111_1101110111, \
	16'b000000_0000011110, \
	16'b111111_1111011111, \
	16'b000000_0001101100, \
	16'b111111_1111111000, \
	16'b000000_0000110101, \
	16'b111111_1101101101, \
	16'b111111_1110000100, \
	16'b000000_0010000011, \
	16'b000000_0000000100, \
	16'b111111_1101011100, \
	16'b111111_1111110111, \
	16'b000000_0000101111, \
	16'b000000_0001000011, \
	16'b000000_0000110101, \
	16'b000000_0000111000, \
	16'b000000_0000000101, \
	16'b000000_0001111001, \
	16'b111111_1111000000, \
	16'b111111_1111101101, \
	16'b000000_0100010100, \
	16'b000000_0001000100, \
	16'b000000_0001100000, \
	16'b000000_0000111101, \
	16'b111111_1111010010, \
	16'b000000_0011110010, \
	16'b000000_0010101001, \
	16'b111111_1111010101, \
	16'b111111_1110111110, \
	16'b000000_0000110011, \
	16'b111111_1111100110, \
	16'b000000_0010011101, \
	16'b111111_1101110001, \
	16'b000000_0010101101, \
	16'b000000_0001101100, \
	16'b111111_1111010001, \
	16'b000000_0101000000, \
	16'b111111_1111100110, \
	16'b000000_0000101000, \
	16'b111111_1111010110, \
	16'b111111_1111011110, \
	16'b000000_0011011100, \
	16'b000000_0010101100, \
	16'b111111_1111111010, \
	16'b000000_0010011011, \
	16'b111111_1111110100, \
	16'b111111_1111101111, \
	16'b111111_1111000101, \
	16'b000000_0001011001, \
	16'b111111_1111111111, \
	16'b000000_0000111101, \
	16'b111111_1100100111, \
	16'b111111_1111111100, \
	16'b000000_0010010111, \
	16'b111111_1111100011, \
	16'b111111_1100100110, \
	16'b000000_0010101110, \
	16'b000000_0010000011, \
	16'b000000_0000001100, \
	16'b111111_1010100110, \
	16'b000000_0001000001, \
	16'b111111_1111110010, \
	16'b111111_1110101101, \
	16'b000000_0001011001, \
	16'b000000_0000101110, \
	16'b000000_0001111100, \
	16'b000000_0010101000, \
	16'b111111_1101011111, \
	16'b000000_0001110111, \
	16'b111111_1101111111, \
	16'b000000_0001100001, \
	16'b000000_0001111000, \
	16'b111111_1010001100, \
	16'b000000_0011110000, \
	16'b000000_0010110001, \
	16'b111111_1111101001, \
	16'b111111_1110101101, \
	16'b111111_1111001110, \
	16'b111111_1111101011, \
	16'b111111_1110111110, \
	16'b111111_1110100000, \
	16'b000000_0001111110, \
	16'b000000_0001010110, \
	16'b111111_1111010100, \
	16'b000000_0010010101, \
	16'b111111_1110101111, \
	16'b000000_0000101101, \
	16'b000000_0000010101, \
	16'b000000_0001010101, \
	16'b000000_0100101101, \
	16'b000000_0010011111, \
	16'b111111_1110110010, \
	16'b000000_0000111010, \
	16'b000000_0000111101, \
	16'b111111_1111100110, \
	16'b000000_0001101010, \
	16'b000000_0011001110, \
	16'b000000_0000100001, \
	16'b000000_0000011101, \
	16'b000000_0010000011, \
	16'b000000_0000001010, \
	16'b000000_0010011010, \
	16'b000000_0000100110, \
	16'b111111_1010110110, \
	16'b000000_0011011010, \
	16'b111111_1111110101, \
	16'b000000_0001000011, \
	16'b111111_1101101000, \
	16'b000000_0001111000, \
	16'b000000_0000010011, \
	16'b111111_1111010100, \
	16'b111111_1100011011, \
	16'b000000_0000110110, \
	16'b000000_0001110010, \
	16'b000000_0011001011, \
	16'b111111_1110100011, \
	16'b000000_0001000010, \
	16'b111111_1000111000, \
	16'b111111_1110100100, \
	16'b111111_1101000000, \
	16'b111111_1001111100, \
	16'b000000_0010111110, \
	16'b000000_0010111111, \
	16'b111111_1111100101, \
	16'b000000_0010111101, \
	16'b111111_1111101111, \
	16'b000000_0000010111, \
	16'b111111_1111111011, \
	16'b111111_1111010110, \
	16'b000000_0001011110, \
	16'b111111_1111111110, \
	16'b111111_1111100100, \
	16'b000000_0000010100, \
	16'b000000_0001110110, \
	16'b000000_0010001111, \
	16'b000000_0000000100, \
	16'b000000_0100100000, \
	16'b000000_0011001011, \
	16'b000000_0000100110, \
	16'b000000_0000110110, \
	16'b111111_1111000111, \
	16'b111111_1110010011, \
	16'b111111_1110011010, \
	16'b111111_1111100100, \
	16'b000000_0100001100, \
	16'b111111_1110000000, \
	16'b111111_1101111111, \
	16'b000000_0100011011, \
	16'b000000_0000000101, \
	16'b000000_0010111011, \
	16'b111111_1111000110, \
	16'b111111_1100110000, \
	16'b000000_0011001111, \
	16'b111111_1011110001, \
	16'b111111_1111100100, \
	16'b000000_0100100111, \
	16'b000000_0000100011, \
	16'b111111_1111110010, \
	16'b000000_0000011000, \
	16'b111111_1011100100, \
	16'b000000_0000101001, \
	16'b111111_1110001011, \
	16'b000000_0000110110, \
	16'b000000_0001011000, \
	16'b000000_0001001011, \
	16'b111111_1010000000, \
	16'b000000_0001111100, \
	16'b111111_1010110000, \
	16'b111111_1111000101, \
	16'b111111_1111101001, \
	16'b000000_0001001101, \
	16'b000000_0000000001, \
	16'b111111_1110110010, \
	16'b111111_1110111110, \
	16'b111111_1111101100, \
	16'b111111_1110101101, \
	16'b000000_0010110011, \
	16'b111111_1111110101, \
	16'b000000_0000101011, \
	16'b111111_1111101110, \
	16'b111111_1110000111, \
	16'b000000_0000101101, \
	16'b111111_1111010101, \
	16'b111111_1110001010, \
	16'b111111_1110001111, \
	16'b000000_0000000110, \
	16'b111111_1101100000, \
	16'b000000_0000111011, \
	16'b111111_1000101100, \
	16'b111111_1111111100, \
	16'b111111_1111111101, \
	16'b111111_1111110010, \
	16'b111111_1010100100, \
	16'b111111_1010001110, \
	16'b111111_1100001011, \
	16'b000000_0100001001, \
	16'b000000_0000111011, \
	16'b000000_1000011111, \
	16'b000000_0000100011, \
	16'b111111_1101001001, \
	16'b000000_0001010100, \
	16'b111111_1011100101, \
	16'b000000_0010000010, \
	16'b000000_0011111100, \
	16'b000000_0000011001, \
	16'b000000_0001000110, \
	16'b111111_1110111101, \
	16'b111111_1011100011, \
	16'b111111_1101111111, \
	16'b111111_1100001101, \
	16'b000000_0000111110, \
	16'b000000_0000010100, \
	16'b111111_1110001110, \
	16'b111111_1000011011, \
	16'b111111_1111010010, \
	16'b111111_1101100011, \
	16'b111111_1011100111, \
	16'b111111_1010111100, \
	16'b111111_1011100001, \
	16'b111111_1111010100, \
	16'b000000_0000111101, \
	16'b000000_0000111100, \
	16'b111111_1110100001, \
	16'b000000_0000101011, \
	16'b000000_0001001110, \
	16'b111111_1110010111, \
	16'b000000_0001010001, \
	16'b111111_1111110001, \
	16'b111111_1111100111, \
	16'b111111_1111000001, \
	16'b000000_0001011011, \
	16'b111111_1111001010, \
	16'b111111_1101101001, \
	16'b000000_0000110010, \
	16'b000000_0000110011, \
	16'b111111_1111101110, \
	16'b111111_1101111010, \
	16'b000000_0001000000, \
	16'b000000_0010010110, \
	16'b111111_1111000001, \
	16'b111111_1110110110, \
	16'b111111_1110001001, \
	16'b111111_1111001011, \
	16'b000000_0000111100, \
	16'b000000_0001100111, \
	16'b000000_0001101110, \
	16'b000000_0010101101, \
	16'b111111_1111010001, \
	16'b000000_0000110010, \
	16'b111111_1111011101, \
	16'b000000_0101100111, \
	16'b000000_0000111111, \
	16'b000000_0001000010, \
	16'b111111_1101110001, \
	16'b000000_0001110000, \
	16'b000000_0000101001, \
	16'b111111_1110000111, \
	16'b000000_0011100111, \
	16'b111111_1111101000, \
	16'b111111_1110010100, \
	16'b111111_1100000001, \
	16'b000000_0000010000, \
	16'b111111_1111111101, \
	16'b111111_1111110110, \
	16'b111111_1010000111, \
	16'b111111_1011111110, \
	16'b111111_1110111100, \
	16'b000000_0000101000, \
	16'b000000_0001000010, \
	16'b000000_0000100110, \
	16'b111111_1110011111, \
	16'b111111_1110010110, \
	16'b000000_0010000001, \
	16'b000000_0000010001, \
	16'b000000_0001111101, \
	16'b000000_0000001001, \
	16'b111111_1110011101, \
	16'b000000_0000001110, \
	16'b000000_0000001011, \
	16'b111111_1111111000, \
	16'b111111_1110011010, \
	16'b000000_0001001111, \
	16'b000000_0000111011, \
	16'b111111_1111110001, \
	16'b111111_1100001001, \
	16'b111111_1111110010, \
	16'b000000_0000000101, \
	16'b111111_1111111100, \
	16'b111111_1110001101, \
	16'b111111_1101101001, \
	16'b111111_1011001101, \
	16'b000000_0000100101, \
	16'b111111_1111111001, \
	16'b000000_0000111100, \
	16'b000000_0001010100, \
	16'b111111_1100111011, \
	16'b000000_0001100010, \
	16'b111111_1110111100, \
	16'b111111_1101011111, \
	16'b000000_0000010111, \
	16'b000000_0000000010, \
	16'b000000_0001110111, \
	16'b111111_1110011000, \
	16'b111111_1110111001, \
	16'b000000_0010110100, \
	16'b000000_0000111000, \
	16'b111111_1111001010, \
	16'b000000_0000100011, \
	16'b000000_0001100000, \
	16'b000000_0010001111, \
	16'b111111_1111100111, \
	16'b000000_0000011101, \
	16'b000000_0001001001, \
	16'b000000_0001001000, \
	16'b111111_1111100100, \
	16'b111111_1111110010, \
	16'b111111_1110100010, \
	16'b000000_0000110110, \
	16'b000000_0000110110, \
	16'b000000_0001101001, \
	16'b000000_0000100001, \
	16'b000000_0000110101, \
	16'b111111_1111110100, \
	16'b111111_1111001100, \
	16'b111111_1111010110, \
	16'b111111_1110010110, \
	16'b111111_1110100111, \
	16'b111111_1110010010, \
	16'b000000_0000111000, \
	16'b111111_1101110000, \
	16'b000000_0001011010, \
	16'b000000_0000011011, \
	16'b000000_0000110000, \
	16'b000000_0001111100, \
	16'b111111_1111011101, \
	16'b111111_1111111101, \
	16'b111111_1101011011, \
	16'b111111_1111101100, \
	16'b111111_1110111101, \
	16'b000000_0010010011, \
	16'b111111_1111010100, \
	16'b000000_0001000001, \
	16'b111111_1110011101, \
	16'b111111_1111110010, \
	16'b000000_0100010010, \
	16'b111111_1111010010, \
	16'b111111_1101011111, \
	16'b000000_0001101100, \
	16'b000000_0000011000, \
	16'b000000_0001000110, \
	16'b000000_0000111010, \
	16'b111111_1110111001, \
	16'b000000_0101001011, \
	16'b111111_1110100001, \
	16'b111111_1011001011, \
	16'b000000_0011001110, \
	16'b111111_1110000011, \
	16'b000000_0010101101, \
	16'b111111_1111110110, \
	16'b000000_0001010110, \
	16'b000000_0111110010, \
	16'b111111_1110011011, \
	16'b111111_1100111101, \
	16'b111111_1111111010, \
	16'b111111_1011011100, \
	16'b111111_1111100001, \
	16'b111111_1111010111, \
	16'b111111_1111100000, \
	16'b000000_0000000010, \
	16'b111111_1100100100, \
	16'b111111_1111000010, \
	16'b111111_1111100011, \
	16'b000000_0000101111, \
	16'b111111_1110110001, \
	16'b111111_1111010111, \
	16'b111111_1111000110, \
	16'b000000_0001011011, \
	16'b111111_1101110101, \
	16'b000000_0000000111, \
	16'b000000_0000100110, \
	16'b111111_1111110011, \
	16'b111111_1111101010, \
	16'b000000_0000111001, \
	16'b000000_0000010110, \
	16'b000000_0011101011, \
	16'b000000_0001010100, \
	16'b000000_0000000001, \
	16'b000000_0001101111, \
	16'b111111_1111000001, \
	16'b000000_0001011001, \
	16'b111111_1110111000, \
	16'b000000_0001110010, \
	16'b000000_0011111010, \
	16'b111111_1111110011, \
	16'b111111_1110001011, \
	16'b000000_0001000001, \
	16'b111111_1111010001, \
	16'b000000_0010110011, \
	16'b111111_1110010101, \
	16'b000000_0010111010, \
	16'b000000_0100001000, \
	16'b111111_1110100001, \
	16'b111111_1011101011, \
	16'b000000_0001011111, \
	16'b111111_1110010010, \
	16'b000000_0100010101, \
	16'b111111_1110111010, \
	16'b000000_0010001000, \
	16'b000000_1000001011, \
	16'b111111_1111000010, \
	16'b111111_1011001010, \
	16'b000000_0000001100, \
	16'b111111_1100101011, \
	16'b111111_1111001000, \
	16'b111111_1111111011, \
	16'b000000_0001101001, \
	16'b000000_0000010000, \
	16'b111111_1011011111, \
	16'b111111_1111111010, \
	16'b111111_1111011001, \
	16'b111111_1111010111, \
	16'b111111_1100010011, \
	16'b111111_1111000011, \
	16'b000000_0000011110, \
	16'b000000_0000100111, \
	16'b111111_1111000111, \
	16'b111111_1110001111, \
	16'b000000_0001001000, \
	16'b111111_1100100100, \
	16'b000000_0010110001, \
	16'b111111_1110111100, \
	16'b000000_0001001110, \
	16'b000000_0011100111, \
	16'b000000_0000000011, \
	16'b111111_1110101000, \
	16'b111111_1111000111, \
	16'b111111_1110000111, \
	16'b000000_0100011101, \
	16'b000000_0001111011, \
	16'b000000_0011010100, \
	16'b000000_0011010101, \
	16'b111111_1111001001, \
	16'b111111_1110001001, \
	16'b111111_1010110000, \
	16'b111111_1111101010, \
	16'b000000_0011000110, \
	16'b000000_0000010101, \
	16'b000000_0001110010, \
	16'b000000_0001111000, \
	16'b111111_1111010011, \
	16'b000000_0001111110, \
	16'b111111_1110001011, \
	16'b000000_0001000111, \
	16'b000000_0010001111, \
	16'b111111_1111111101, \
	16'b000000_0010001111, \
	16'b111111_1101110101, \
	16'b000000_0000111111, \
	16'b111111_1111001011, \
	16'b111111_1110111110, \
	16'b000000_0000011011, \
	16'b111111_1111110100, \
	16'b000000_0000101010, \
	16'b000000_0001100101, \
	16'b111111_1111001100, \
	16'b000000_0000000100, \
	16'b111111_1111001010, \
	16'b111111_1111111001, \
	16'b111111_1011001100, \
	16'b111111_1110111110, \
	16'b111111_1110010010, \
	16'b111111_1110011011, \
	16'b111111_1100101000, \
	16'b111111_1111000111, \
	16'b111111_1010100010, \
	16'b000000_0001110011, \
	16'b111111_1100011011, \
	16'b000000_1011010011, \
	16'b111111_1111010101, \
	16'b111111_1111110110, \
	16'b000000_0011011110, \
	16'b111111_1101001111, \
	16'b111111_1101110111, \
	16'b111111_1110000011, \
	16'b000000_0000000011, \
	16'b000000_0101100101, \
	16'b111111_1110011000, \
	16'b000000_0001000011, \
	16'b000000_0010001000, \
	16'b111111_1110001110, \
	16'b111111_1101100010, \
	16'b111111_1011100000, \
	16'b000000_0000101000, \
	16'b000000_0001110011, \
	16'b111111_1110101010, \
	16'b111111_1101110010, \
	16'b000000_0000001001, \
	16'b111111_1111101000, \
	16'b111111_1111101110, \
	16'b111111_1110100111, \
	16'b000000_0001010101, \
	16'b111111_1110001110, \
	16'b000000_0000111000, \
	16'b000000_0001100011, \
	16'b000000_0000010111, \
	16'b000000_0011110110, \
	16'b000000_0001101010, \
	16'b111111_1110111000, \
	16'b000000_0001000010, \
	16'b111111_1110111010, \
	16'b000000_0000010011, \
	16'b000000_0000111111, \
	16'b000000_0001000000, \
	16'b000000_0001100010, \
	16'b000000_0001110100, \
	16'b111111_1111010001, \
	16'b000000_0001001010, \
	16'b111111_1111001110, \
	16'b000000_0001101011, \
	16'b111111_1110110110, \
	16'b111111_1100111110, \
	16'b000000_0001010100, \
	16'b000000_0000000011, \
	16'b111111_1111111111, \
	16'b000000_0001101001, \
	16'b000000_0110010100, \
	16'b000000_0000011001, \
	16'b000000_0000000000, \
	16'b000000_0010101000, \
	16'b000000_0001010110, \
	16'b000000_0010011110, \
	16'b111111_1111100110, \
	16'b000000_0000001110, \
	16'b000000_0100111011, \
	16'b111111_1111001011, \
	16'b000000_0000001000, \
	16'b000000_0000000010, \
	16'b111111_1101110111, \
	16'b111111_1100111101, \
	16'b111111_1101100010, \
	16'b000000_0000001110, \
	16'b111111_1011010110, \
	16'b000000_0000010010, \
	16'b111111_1111101010, \
	16'b000000_0000001010, \
	16'b111111_1101011010, \
	16'b111111_1110100010, \
	16'b111111_1111101101, \
	16'b000000_0011110001, \
	16'b111111_1101111011, \
	16'b111111_1111001101, \
	16'b111111_1110010100, \
	16'b000000_0001101010, \
	16'b000000_0100010100, \
	16'b000000_0010011111, \
	16'b000000_0000100010, \
	16'b000000_0001110110, \
	16'b000000_0001000101, \
	16'b111111_1110101010, \
	16'b000000_0001000100, \
	16'b000000_0000001010, \
	16'b111111_1111100001, \
	16'b111111_1101110110, \
	16'b000000_0000001111, \
	16'b000000_0000001000, \
	16'b111111_1110010011, \
	16'b111111_1111001001, \
	16'b000000_0000101000, \
	16'b000000_0000101100, \
	16'b111111_1101100110, \
	16'b111111_1101011101, \
	16'b000000_0000000000, \
	16'b111111_1111000001, \
	16'b111111_1110011001, \
	16'b000000_0000011111, \
	16'b111111_1110011011, \
	16'b000000_0001000110, \
	16'b111111_1011101100, \
	16'b111111_1111011001, \
	16'b000000_0000011111, \
	16'b000000_0011000011, \
	16'b000000_0001001110, \
	16'b000000_0000000000, \
	16'b000000_0011101100, \
	16'b111111_1101101010, \
	16'b000000_0000111011, \
	16'b000000_0011100001, \
	16'b000000_0000110011, \
	16'b111111_1111110010, \
	16'b111111_1110010001, \
	16'b000000_0000001101, \
	16'b000000_0011110110, \
	16'b000000_0000010100, \
	16'b111111_1111110101, \
	16'b000000_0000001001, \
	16'b000000_0000001111, \
	16'b111111_1100010000, \
	16'b111111_1010100010, \
	16'b111111_1110110111, \
	16'b111111_1110011011, \
	16'b111111_1101110100, \
	16'b111111_1011000111, \
	16'b111111_1101100110, \
	16'b111111_1111000111, \
	16'b000000_0000011000, \
	16'b000000_0000001101, \
	16'b000000_0001101011, \
	16'b000000_0010011011, \
	16'b111111_1110101000, \
	16'b111111_1101110011, \
	16'b111111_1110110000, \
	16'b111111_1111110010, \
	16'b111111_1110111100, \
	16'b111111_1111100111, \
	16'b111111_1111110111, \
	16'b000000_0000000000, \
	16'b000000_0000001101, \
	16'b000000_0000100101, \
	16'b111111_1101010100, \
	16'b000000_0001010000, \
	16'b111111_1011000010, \
	16'b000000_0010000001, \
	16'b111111_1101001101, \
	16'b000000_0001000111, \
	16'b000000_0000011101, \
	16'b111111_1101100000, \
	16'b111111_1101011001, \
	16'b111111_1111101000, \
	16'b111111_1101111110, \
	16'b111111_1111100011, \
	16'b000000_0001000110, \
	16'b000000_0001011011, \
	16'b111111_1010010100, \
	16'b000000_0000011001, \
	16'b000000_0001100000, \
	16'b000000_0000001101, \
	16'b111111_1100111010, \
	16'b111111_1110011100, \
	16'b000000_0001111000, \
	16'b111111_1111101001, \
	16'b111111_1000110001, \
	16'b000000_0000000100, \
	16'b111111_1100111010, \
	16'b111111_1110001000, \
	16'b000000_0000001011, \
	16'b000000_0001111101, \
	16'b000000_0000000100, \
	16'b111111_1110100011, \
	16'b111111_1111101010, \
	16'b000000_0000011000, \
	16'b000000_0000011000, \
	16'b111111_1111111011, \
	16'b000000_0000110101, \
	16'b000000_0011110010, \
	16'b000000_0000111101, \
	16'b000000_0010010000, \
	16'b000000_0000110101, \
	16'b000000_0010000100, \
	16'b111111_1111010000, \
	16'b000000_0000010111, \
	16'b000000_0010110100, \
	16'b000000_0011010110, \
	16'b111111_1111101011, \
	16'b000000_0000000011, \
	16'b000000_0010000010, \
	16'b000000_0011001001, \
	16'b000000_0001001011, \
	16'b000000_0010000000, \
	16'b000000_0001010111, \
	16'b000000_0111100111, \
	16'b111111_1110100101, \
	16'b111111_1111001111, \
	16'b000000_0111101000, \
	16'b000000_0010001101, \
	16'b111111_1111110000, \
	16'b111111_1101111110, \
	16'b000000_0000100001, \
	16'b000000_0010110000, \
	16'b111111_1110111011, \
	16'b111111_1100110110, \
	16'b000000_0001110110, \
	16'b000000_0000001010, \
	16'b000000_0000000000, \
	16'b111111_1100011101, \
	16'b000000_0001001010, \
	16'b000000_0001100110, \
	16'b111111_1101111000, \
	16'b111111_1101010000, \
	16'b111111_1001001100, \
	16'b000000_0010001110, \
	16'b111111_1111111001, \
	16'b111111_1101111011, \
	16'b000000_0100110100, \
	16'b000000_0010000011, \
	16'b111111_1110010001, \
	16'b111111_1110011111, \
	16'b111111_1011110011, \
	16'b000000_0010110000, \
	16'b000000_0100110100, \
	16'b000000_0001010011, \
	16'b000000_0010000011, \
	16'b000000_0010001110, \
	16'b000000_0000100101, \
	16'b000000_0000010000, \
	16'b111111_1111111110, \
	16'b000000_0011001111, \
	16'b111111_1111101000, \
	16'b111111_1111110011, \
	16'b000000_0001101001, \
	16'b000000_0011010100, \
	16'b111111_1111101100, \
	16'b000000_0000111101, \
	16'b000000_0011011001, \
	16'b000000_0000101110, \
	16'b000000_0010011001, \
	16'b111111_1111101000, \
	16'b000000_0100010110, \
	16'b000000_0101011100, \
	16'b000000_0000010101, \
	16'b111111_1110001100, \
	16'b000000_0010101100, \
	16'b000000_0010100100, \
	16'b000000_0001101000, \
	16'b111111_1100110100, \
	16'b000000_0010000001, \
	16'b111111_1101101110, \
	16'b111111_1111010110, \
	16'b000000_0001111001, \
	16'b000000_0000001110, \
	16'b111111_1111010000, \
	16'b000000_0001100111, \
	16'b111111_0111100011, \
	16'b000000_0001100000, \
	16'b111111_1011101001, \
	16'b000000_0100001000, \
	16'b111111_1010111101, \
	16'b111111_1101010111, \
	16'b000000_0001001010, \
	16'b000000_0011000100, \
	16'b000000_0001010001, \
	16'b000000_0100001000, \
	16'b111111_1110110111, \
	16'b111111_1110110000, \
	16'b111111_1110001101, \
	16'b111111_1101111110, \
	16'b000000_0010101010, \
	16'b000000_0001000100, \
	16'b000000_0000100001, \
	16'b111111_1101001011, \
	16'b000000_0000010110, \
	16'b000000_0000111100, \
	16'b000000_0000101101, \
	16'b000000_0000011101, \
	16'b000000_0000010000, \
	16'b000000_0000110001, \
	16'b000000_0000010010, \
	16'b111111_1101101101, \
	16'b000000_0000000100, \
	16'b000000_0000111000, \
	16'b111111_1111010011, \
	16'b111111_1101110100, \
	16'b111111_1110100011, \
	16'b000000_0000010101, \
	16'b000000_0000000101, \
	16'b111111_1111110101, \
	16'b111111_1100010001, \
	16'b111111_1111000011, \
	16'b111111_1111100001, \
	16'b000000_0000001010, \
	16'b111111_1101010010, \
	16'b111111_1111100111, \
	16'b000000_0000101100, \
	16'b000000_0000001110, \
	16'b111111_0100011101, \
	16'b000000_0000101001, \
	16'b111111_1110111100, \
	16'b111111_1111010010, \
	16'b111111_1110011000, \
	16'b000000_0001110100, \
	16'b000000_0000111010, \
	16'b111111_1111110100, \
	16'b111111_0101001000, \
	16'b000000_0101110111, \
	16'b111111_1110101111, \
	16'b111111_1110001001, \
	16'b000000_0000000010, \
	16'b000000_0101011000, \
	16'b111111_1111101110, \
	16'b000000_0001010010, \
	16'b111111_1000001110, \
	16'b000000_0001000110, \
	16'b111111_1101011001, \
	16'b111111_1101001111, \
	16'b000000_0100000111, \
	16'b000000_0001101000, \
	16'b111111_1111010011, \
	16'b111111_1111110000, \
	16'b111111_1110010100, \
	16'b111111_1110110010, \
	16'b111111_1101111110, \
	16'b111111_1111011001, \
	16'b111111_1110101101, \
	16'b111111_1111100100, \
	16'b111111_1111001110, \
	16'b111111_1111100000, \
	16'b111111_1110110000, \
	16'b000000_0001110101, \
	16'b111111_1110000110, \
	16'b000000_0000100101, \
	16'b111111_1110111111, \
	16'b111111_1110111100, \
	16'b000000_0000001001, \
	16'b111111_1110101011, \
	16'b111111_1111110000, \
	16'b111111_1111000010, \
	16'b000000_0001011110, \
	16'b111111_1100010001, \
	16'b111111_1110101111, \
	16'b111111_1101001001, \
	16'b000000_0001011101, \
	16'b111111_1110000010, \
	16'b111111_1110110000, \
	16'b000000_0000011111, \
	16'b111111_1111001011, \
	16'b111111_1111000010, \
	16'b111111_1100001110, \
	16'b000000_0010111101, \
	16'b111111_1111111111, \
	16'b000000_0000010111, \
	16'b111111_1101111010, \
	16'b000000_0010101000, \
	16'b111111_1111001000, \
	16'b111111_1110101101, \
	16'b000000_0010011000, \
	16'b000000_0101000111, \
	16'b000000_0000011010, \
	16'b000000_0000100110, \
	16'b111111_1101101100, \
	16'b000000_0000000111, \
	16'b111111_1101111101, \
	16'b000000_0000110010, \
	16'b000000_0010111010, \
	16'b000000_0010110111, \
	16'b000000_0000101101, \
	16'b111111_1101111010, \
	16'b000000_0001111110, \
	16'b000000_0001111110, \
	16'b000000_0000101101, \
	16'b000000_0001111111, \
	16'b000000_0000100001, \
	16'b000000_0001001111, \
	16'b111111_1111010010, \
	16'b111111_1110110111, \
	16'b111111_1101100100, \
	16'b111111_1101011010, \
	16'b111111_1110011101, \
	16'b111111_1110110000, \
	16'b111111_1101100101, \
	16'b000000_0000000110, \
	16'b111111_1110011101, \
	16'b111111_1110001010, \
	16'b000000_0000000111, \
	16'b000000_0000000010, \
	16'b111111_1110110010, \
	16'b111111_1101010000, \
	16'b111111_1101010000, \
	16'b111111_1101100111, \
	16'b111111_1111100111, \
	16'b000000_0000110111, \
	16'b000000_0001010111, \
	16'b111111_1110100000, \
	16'b111111_1100001000, \
	16'b111111_1111010001, \
	16'b111111_1110111001, \
	16'b111111_1111110101, \
	16'b111111_1110111100, \
	16'b000000_0000001100, \
	16'b000000_0010100000, \
	16'b111111_1111000001, \
	16'b000000_0001000010, \
	16'b000000_0111000100, \
	16'b000000_0010000101, \
	16'b111111_1111001001, \
	16'b111111_1111110001, \
	16'b111111_1111110000, \
	16'b000000_0011000110, \
	16'b111111_1111111111, \
	16'b000000_0000110100, \
	16'b000000_0000011110, \
	16'b000000_0010010110, \
	16'b111111_1110010011, \
	16'b111111_1110110100, \
	16'b000000_0000100000, \
	16'b111111_1101110111, \
	16'b111111_1110001111, \
	16'b111111_1111010100, \
	16'b000000_0000010110, \
	16'b111111_1110110101, \
	16'b111111_1111001101, \
	16'b111111_1101111000, \
	16'b111111_1110010011, \
	16'b000000_0000000111, \
	16'b111111_1101011100, \
	16'b111111_1111110000, \
	16'b000000_0001100100, \
	16'b111111_1101011111, \
	16'b111111_1101110011, \
	16'b111111_1101111000, \
	16'b000000_0001000110, \
	16'b000000_0000011000, \
	16'b111111_1110001100, \
	16'b111111_1110001001, \
	16'b111111_1110111010, \
	16'b111111_1111011111, \
	16'b000000_0000011011, \
	16'b111111_1111111011, \
	16'b000000_0000011011, \
	16'b000000_0001100110, \
	16'b111111_1110111111, \
	16'b111111_1011001001, \
	16'b000000_0011111010, \
	16'b000000_0001001001, \
	16'b111111_1111011000, \
	16'b000000_0000111100, \
	16'b000000_0001010000, \
	16'b000000_0001111101, \
	16'b111111_1110101010, \
	16'b000000_0000100011, \
	16'b000000_0110100011, \
	16'b111111_1111000010, \
	16'b111111_1101000100, \
	16'b000000_0001101111, \
	16'b111111_1111000101, \
	16'b000000_0010001010, \
	16'b111111_1111101101, \
	16'b000000_0001001101, \
	16'b000000_0110101100, \
	16'b111111_1110010000, \
	16'b111111_1111111011, \
	16'b111111_1110111011, \
	16'b111111_1110101001, \
	16'b000000_0010011100, \
	16'b111111_1110110111, \
	16'b111111_1111001010, \
	16'b000000_0010101111, \
	16'b111111_1110101001, \
	16'b000000_0001100011, \
	16'b111111_1110001000, \
	16'b000000_0001000010, \
	16'b111111_1111110100, \
	16'b000000_0000000101, \
	16'b111111_1101010100, \
	16'b111111_1111000100, \
	16'b111111_1111111011, \
	16'b111111_1110000110, \
	16'b111111_1111011111, \
	16'b111111_1110110101, \
	16'b111111_1110110011, \
	16'b111111_1111101010, \
	16'b111111_1110111100, \
	16'b000000_0001000101, \
	16'b000000_0000101011, \
	16'b111111_1111101000, \
	16'b111111_1011101010, \
	16'b111111_1111111010, \
	16'b000000_0000101101, \
	16'b111111_1101001100, \
	16'b000000_0001101010, \
	16'b000000_0001111000, \
	16'b000000_0000101100, \
	16'b111111_1110110110, \
	16'b111111_1110011100, \
	16'b000000_0000000111, \
	16'b000000_0011101011, \
	16'b111111_1101011100, \
	16'b000000_0100110000, \
	16'b000000_0100100100, \
	16'b000000_0001101010, \
	16'b111111_1001101101, \
	16'b000000_0001110110, \
	16'b111111_1011001111, \
	16'b000000_0100000001, \
	16'b111111_1111000010, \
	16'b000000_0011001110, \
	16'b000000_0100101100, \
	16'b111111_1101000111, \
	16'b111111_1101010011, \
	16'b111111_1110111001, \
	16'b111111_1110110000, \
	16'b111111_1110001110, \
	16'b111111_1101100000, \
	16'b111111_1110101011, \
	16'b000000_0000110011, \
	16'b111111_1101000100, \
	16'b000000_0000000101, \
	16'b111111_1110010010, \
	16'b111111_1111100110, \
	16'b000000_0001000011, \
	16'b000000_0000001000, \
	16'b111111_1101101111, \
	16'b111111_1111001111, \
	16'b000000_0001010011, \
	16'b111111_1111101110, \
	16'b111111_1110001011, \
	16'b000000_0000100110, \
	16'b000000_0000000001, \
	16'b111111_1111110000, \
	16'b111111_1110110010, \
	16'b111111_1110111000, \
	16'b111111_1110001100, \
	16'b000000_0000101010, \
	16'b111111_1101010101, \
	16'b000000_0001010000, \
	16'b000000_0000111101, \
	16'b111111_1111011001, \
	16'b111111_1011111100, \
	16'b000000_0000010000, \
	16'b000000_0000011010, \
	16'b000000_0000001000, \
	16'b000000_0100000100, \
	16'b000000_0000110010, \
	16'b000000_0011000111, \
	16'b111111_1100111011, \
	16'b000000_0000101101, \
	16'b000000_0100110100, \
	16'b111111_1111010111, \
	16'b111111_0110010010, \
	16'b000000_0010011111, \
	16'b111111_1001100101, \
	16'b000000_0100110100, \
	16'b000000_0000100010, \
	16'b000000_0010000110, \
	16'b000000_0101111111, \
	16'b111111_1010101110, \
	16'b111111_1010000001, \
	16'b111111_1101101011, \
	16'b111111_1011111100, \
	16'b111111_1101111011, \
	16'b000000_0000001111, \
	16'b111111_1110010111, \
	16'b111111_1101100110, \
	16'b111111_1011010100, \
	16'b000000_0000011000, \
	16'b111111_1110101100, \
	16'b111111_1111111110, \
	16'b000000_0000110101, \
	16'b111111_1111000110, \
	16'b000000_0000000000, \
	16'b111111_1111011011, \
	16'b111111_1111011010, \
	16'b000000_0000011011, \
	16'b111111_1101011010, \
	16'b000000_0001101001, \
	16'b111111_1101101110, \
	16'b000000_0000100100, \
	16'b111111_1101010111, \
	16'b111111_1111011011, \
	16'b000000_0001011101, \
	16'b000000_0000101101, \
	16'b111111_1101110011, \
	16'b000000_0001100000, \
	16'b000000_0010001010, \
	16'b000000_0001100111, \
	16'b111111_1100101101, \
	16'b000000_0000010111, \
	16'b000000_0001001111, \
	16'b000000_0000111110, \
	16'b000000_0001001100, \
	16'b111111_1111001000, \
	16'b000000_0100010011, \
	16'b111111_1110010001, \
	16'b000000_0100000100, \
	16'b000000_0001010001, \
	16'b000000_0000111111, \
	16'b111111_1001001000, \
	16'b000000_0000001000, \
	16'b111111_1100111000, \
	16'b000000_0101100010, \
	16'b111111_1111100011, \
	16'b000000_0101110000, \
	16'b000000_0000110111, \
	16'b111111_1101000100, \
	16'b111111_1000101110, \
	16'b111111_1101101000, \
	16'b111111_1101101101, \
	16'b000000_0000001010, \
	16'b000000_0000101110, \
	16'b111111_1111111010, \
	16'b000000_0001100001, \
	16'b111111_1101010000, \
	16'b000000_0001100001, \
	16'b111111_1101111101, \
	16'b000000_0000010010, \
	16'b000000_0010001000, \
	16'b111111_1110100110, \
	16'b111111_1111011111, \
	16'b000000_0001000011, \
	16'b000000_0000100010, \
	16'b111111_1101110100, \
	16'b111111_1110010110, \
	16'b000000_0000101001, \
	16'b111111_1100011111, \
	16'b111111_1111100111, \
	16'b111111_1111100010, \
	16'b000000_0001100111, \
	16'b000000_0000100010, \
	16'b000000_0001110010, \
	16'b111111_1110100010, \
	16'b000000_0001000001, \
	16'b111111_1111111010, \
	16'b111111_1110010001, \
	16'b111111_1101110110, \
	16'b000000_0000001000, \
	16'b000000_0010110001, \
	16'b000000_0010001111, \
	16'b111111_1110110111, \
	16'b000000_0001110001, \
	16'b000000_0100010001, \
	16'b111111_1111111101, \
	16'b000000_0001010100, \
	16'b000000_0001101001, \
	16'b000000_0010010100, \
	16'b000000_0000111010, \
	16'b111111_1111101001, \
	16'b111111_1110010000, \
	16'b000000_0011001000, \
	16'b111111_1111111010, \
	16'b000000_0010110011, \
	16'b000000_0000011011, \
	16'b000000_0001010100, \
	16'b111111_1100100011, \
	16'b111111_1110101000, \
	16'b111111_1111010001, \
	16'b000000_0001110010, \
	16'b111111_1111000111, \
	16'b000000_0000011001, \
	16'b111111_1111100100, \
	16'b111111_1111001000, \
	16'b000000_0001100011, \
	16'b000000_0000110010, \
	16'b000000_0001110100, \
	16'b000000_0000100101, \
	16'b000000_0001100110, \
	16'b111111_1111101110, \
	16'b000000_0011010110, \
	16'b000000_0011001001, \
	16'b000000_0011000110, \
	16'b111111_1111000111, \
	16'b000000_0000001110, \
	16'b000000_0011010001, \
	16'b000000_0000001001, \
	16'b111111_1111011010, \
	16'b000000_0111111010, \
	16'b000000_0101000010, \
	16'b111111_1110010110, \
	16'b000000_0000000000, \
	16'b111111_1101010000, \
	16'b000000_0000111010, \
	16'b111111_1110101011, \
	16'b000000_0000100111, \
	16'b111111_1101000111, \
	16'b000000_0000001100, \
	16'b111111_1000110010, \
	16'b000000_0000000011, \
	16'b000000_0000111000, \
	16'b000000_0001001111, \
	16'b111111_1110001010, \
	16'b111111_1100000110, \
	16'b111111_1011101001, \
	16'b111111_1111101111, \
	16'b111111_1111001010, \
	16'b000000_0001010110, \
	16'b000000_0010110110, \
	16'b000000_0001100000, \
	16'b000000_0001111100, \
	16'b000000_0000011000, \
	16'b000000_0010000111, \
	16'b000000_0001100100, \
	16'b000000_0010100101, \
	16'b000000_0000000000, \
	16'b000000_0000010110, \
	16'b111111_1111011001, \
	16'b000000_0001001110, \
	16'b000000_0000010101, \
	16'b111111_1110000001, \
	16'b000000_0000100101, \
	16'b111111_1101111010, \
	16'b000000_0000000011, \
	16'b000000_0000111101, \
	16'b111111_1111111111, \
	16'b111111_1111110101, \
	16'b000000_0001011110, \
	16'b000000_0110101010, \
	16'b111111_1111011001, \
	16'b111111_1111111111, \
	16'b000000_0000100011, \
	16'b000000_0001100000, \
	16'b000000_0100010011, \
	16'b000000_0001001001, \
	16'b000000_0000001111, \
	16'b000000_1001110011, \
	16'b000000_0000110100, \
	16'b111111_1110010100, \
	16'b111111_1110011010, \
	16'b111111_1111011010, \
	16'b000000_0001010011, \
	16'b111111_1101001110, \
	16'b000000_0001001000, \
	16'b000000_0011011001, \
	16'b000000_0000000111, \
	16'b111111_1101100000, \
	16'b000000_0100011010, \
	16'b000000_0011001011, \
	16'b000000_0000100011, \
	16'b111111_1111110001, \
	16'b111111_1011100110, \
	16'b000000_0010011000, \
	16'b000000_0000101100, \
	16'b111111_1101000110, \
	16'b000000_0010111100, \
	16'b000000_0010000000, \
	16'b000000_0010101110, \
	16'b000000_0001100100, \
	16'b000000_0000100100, \
	16'b000000_0011101011, \
	16'b111111_1111110111, \
	16'b111111_1110111101, \
	16'b111111_1111110010, \
	16'b111111_1111111000, \
	16'b111111_1111001001, \
	16'b111111_1111101110, \
	16'b000000_0000001001, \
	16'b111111_1101100111, \
	16'b111111_1101010110, \
	16'b111111_1111000111, \
	16'b111111_1111111010, \
	16'b111111_1101001001, \
	16'b000000_0001000011, \
	16'b111111_1111011100, \
	16'b000000_0001100001, \
	16'b000000_0000110110, \
	16'b111111_1110001000, \
	16'b111111_1110000001, \
	16'b000000_0010101011, \
	16'b111111_1111001101, \
	16'b000000_0011110100, \
	16'b000000_0000100010, \
	16'b111111_1111000101, \
	16'b000000_0011010111, \
	16'b111111_1011110011, \
	16'b111111_1111101010, \
	16'b000000_0100111100, \
	16'b000000_0000011000, \
	16'b000000_0000101000, \
	16'b000000_0011100111, \
	16'b111111_1100001010, \
	16'b000000_0010010110, \
	16'b111111_1100110110, \
	16'b000000_0000100111, \
	16'b000000_0101001000, \
	16'b000000_0000001010, \
	16'b111111_1110111011, \
	16'b000000_0010001000, \
	16'b111111_1011000001, \
	16'b000000_0010011011, \
	16'b111111_1100111110, \
	16'b111111_1100110011, \
	16'b000000_0010110001, \
	16'b111111_1110101101, \
	16'b111111_1110100011, \
	16'b000000_0000100100, \
	16'b111111_1100110010, \
	16'b000000_0101001111, \
	16'b111111_1011011101, \
	16'b111111_1101111111, \
	16'b000000_0000101101, \
	16'b111111_1100111100, \
	16'b111111_1101110110, \
	16'b111111_1111001100, \
	16'b111111_1111100011, \
	16'b000000_0001001010, \
	16'b111111_1110100010, \
	16'b111111_1110001011, \
	16'b111111_1111111011, \
	16'b111111_1100110001, \
	16'b000000_0000000101, \
	16'b111111_1111001010, \
	16'b000000_0000110100, \
	16'b111111_1110011010, \
	16'b111111_1111001100, \
	16'b000000_0000101010, \
	16'b111111_1111110010, \
	16'b111111_1111000101, \
	16'b111111_1110001001, \
	16'b111111_1111000111, \
	16'b000000_0001111111, \
	16'b111111_1110101110, \
	16'b111111_1111000001, \
	16'b000000_0000101001, \
	16'b000000_0100000010, \
	16'b111111_1111110001, \
	16'b000000_0000000000, \
	16'b000000_0011100100, \
	16'b000000_0010011101, \
	16'b000000_0001011001, \
	16'b111111_1111110111, \
	16'b000000_0001000001, \
	16'b000000_0100100110, \
	16'b111111_1101111011, \
	16'b000000_0011000011, \
	16'b111111_1111110010, \
	16'b000000_0001101110, \
	16'b000000_0001001101, \
	16'b111111_1101011111, \
	16'b111111_1110101011, \
	16'b000000_0001110001, \
	16'b111111_1011101010, \
	16'b000000_0010111001, \
	16'b000000_0000000101, \
	16'b000000_0010100000, \
	16'b000000_0001001000, \
	16'b111111_1001110001, \
	16'b111111_1110000101, \
	16'b111111_1111010101, \
	16'b111111_1101111100, \
	16'b000000_0000000011, \
	16'b111111_1110111101, \
	16'b111111_1111101000, \
	16'b111111_1110111111, \
	16'b111111_1110010011, \
	16'b000000_0001000101, \
	16'b000000_0000001110, \
	16'b111111_1110111101, \
	16'b000000_0001001001, \
	16'b000000_0001011010, \
	16'b000000_0000010101, \
	16'b111111_1101111110, \
	16'b000000_0000000001, \
	16'b111111_1101110100, \
	16'b000000_0001001100, \
	16'b111111_1110011100, \
	16'b111111_1001100101, \
	16'b111111_1111111110, \
	16'b000000_0010101110, \
	16'b111111_1110011011, \
	16'b111111_1111100011, \
	16'b111111_1111000101, \
	16'b000000_0001010100, \
	16'b111111_1110011010, \
	16'b000000_0000100010, \
	16'b000000_0001010001, \
	16'b000000_0100000100, \
	16'b000000_0000001011, \
	16'b111111_1111011100, \
	16'b111111_1111111000, \
	16'b000000_0000101100, \
	16'b111111_1111011111, \
	16'b000000_0011000010, \
	16'b111111_1111101111, \
	16'b000000_0010110010, \
	16'b000000_0000001000, \
	16'b111111_1110100001, \
	16'b111111_1101101011, \
	16'b000000_0000101001, \
	16'b111111_1110000100, \
	16'b000000_0100010110, \
	16'b111111_1111111010, \
	16'b000000_0010111011, \
	16'b000000_0000100110, \
	16'b111111_1110010110, \
	16'b111111_1101010101, \
	16'b111111_1111100111, \
	16'b000000_0001011111, \
	16'b000000_0001000111, \
	16'b000000_0000000111, \
	16'b111111_1110101100, \
	16'b000000_0000011000, \
	16'b111111_1111101000, \
	16'b111111_1111000100, \
	16'b000000_0000000000, \
	16'b111111_1101101010, \
	16'b111111_1101111110, \
	16'b111111_1110101011, \
	16'b111111_1111111110, \
	16'b000000_0000101111, \
	16'b111111_1111011001, \
	16'b000000_0000110101, \
	16'b000000_0000001001, \
	16'b111111_1101101110, \
	16'b111111_1111001110, \
	16'b000000_0001011011, \
	16'b000000_0001100100, \
	16'b111111_1111010000, \
	16'b111111_1110101001, \
	16'b111111_1110011100, \
	16'b000000_0000111010, \
	16'b111111_1111010001, \
	16'b111111_1110100011, \
	16'b111111_1111100101, \
	16'b000000_0000111101, \
	16'b111111_1110111000, \
	16'b111111_1110110111, \
	16'b000000_0010001011, \
	16'b000000_0000011001, \
	16'b111111_1111111011, \
	16'b111111_1100010111, \
	16'b000000_0001000110, \
	16'b000000_0001110001, \
	16'b000000_0000010100, \
	16'b111111_1101101010, \
	16'b111111_1100111000, \
	16'b111111_1111111100, \
	16'b111111_1101000101, \
	16'b111111_1110111010, \
	16'b000000_0000010010, \
	16'b000000_0001110001, \
	16'b111111_1110100110, \
	16'b111111_1100000101, \
	16'b111111_1101110010, \
	16'b000000_0000100000, \
	16'b111111_1101110101, \
	16'b000000_0000011011, \
	16'b111111_1111100001, \
	16'b111111_1110111001, \
	16'b111111_1110001000, \
	16'b111111_1101110111, \
	16'b111111_1111100000, \
	16'b000000_0010111101, \
	16'b000000_0000001010, \
	16'b000000_0000111000, \
	16'b000000_0000000100, \
	16'b000000_0000011001, \
	16'b111111_1110010010, \
	16'b111111_1110001000, \
	16'b111111_1110000101, \
	16'b000000_0001010000, \
	16'b111111_1111001000, \
	16'b111111_1101111111, \
	16'b111111_1111111100, \
	16'b000000_0001010001, \
	16'b111111_1111001110, \
	16'b111111_1110101011, \
	16'b000000_0000000000, \
	16'b000000_0011111011, \
	16'b000000_0000011011, \
	16'b111111_1111010010, \
	16'b000000_0010001101, \
	16'b000000_0011011100, \
	16'b000000_0000010100, \
	16'b111111_1111100101, \
	16'b000000_0000011101, \
	16'b000000_0010111101, \
	16'b111111_1101111010, \
	16'b111111_1111001000, \
	16'b000000_0010011011, \
	16'b000000_0001100111, \
	16'b111111_1111111001, \
	16'b111111_1110101101, \
	16'b000000_0000111111, \
	16'b000000_0011010000, \
	16'b000000_0000111010, \
	16'b111111_1110100100, \
	16'b000000_0000001011, \
	16'b111111_1110111100, \
	16'b111111_1111011101, \
	16'b000000_0000010000, \
	16'b111111_1111011101, \
	16'b000000_0000111011, \
	16'b111111_1111110000, \
	16'b000000_0010000001, \
	16'b000000_0010110001, \
	16'b000000_0001100000, \
	16'b111111_1111111110, \
	16'b111111_1111011011, \
	16'b111111_1101111101, \
	16'b000000_0011010100, \
	16'b111111_1110110100, \
	16'b111111_1111000011, \
	16'b000000_0010000111, \
	16'b000000_0000111010, \
	16'b111111_1111001100, \
	16'b000000_0000000010, \
	16'b111111_1110010111, \
	16'b000000_0010111011, \
	16'b111111_1111101110, \
	16'b111111_1011000111, \
	16'b111111_1111111000, \
	16'b000000_0010111011, \
	16'b111111_1011110000, \
	16'b111111_1100011000, \
	16'b111111_1111100110, \
	16'b000000_0100010001, \
	16'b111111_1101100101, \
	16'b111111_1100110100, \
	16'b000000_0001000011, \
	16'b000000_0011001111, \
	16'b111111_1110000100, \
	16'b111111_1110111101, \
	16'b000000_0000110100, \
	16'b000000_0001011011, \
	16'b111111_1111001100, \
	16'b111111_1100010011, \
	16'b000000_0100010111, \
	16'b000000_0011010111, \
	16'b111111_1100010000, \
	16'b111111_1111110101, \
	16'b000000_0000100111, \
	16'b000000_0001000100, \
	16'b111111_1110101111, \
	16'b111111_1100010011, \
	16'b000000_0001010100, \
	16'b111111_1101110111, \
	16'b111111_1111000110, \
	16'b111111_1111001000, \
	16'b000000_0000111011, \
	16'b000000_0001011010, \
	16'b000000_0000011101, \
	16'b111111_1101010011, \
	16'b000000_0010100010, \
	16'b000000_0000110001, \
	16'b000000_0000011100, \
	16'b000000_0000011010, \
	16'b000000_0000011001, \
	16'b000000_0011000100, \
	16'b000000_0000010110, \
	16'b111111_1111000010, \
	16'b111111_1111001110, \
	16'b111111_1111111101, \
	16'b000000_0001011100, \
	16'b111111_1100110110, \
	16'b111111_1111001100, \
	16'b000000_0010100010, \
	16'b111111_1110001001, \
	16'b111111_1101011011, \
	16'b000000_0001101010, \
	16'b000000_0010000001, \
	16'b111111_1010011111, \
	16'b111111_1101011111, \
	16'b111111_1110110101, \
	16'b000000_0010111101, \
	16'b111111_1110001110, \
	16'b111111_1000011001, \
	16'b000000_0010100110, \
	16'b000000_0100001111, \
	16'b111111_1011000100, \
	16'b111111_1101001110, \
	16'b000000_0000100111, \
	16'b000000_0011100011, \
	16'b111111_1110100110, \
	16'b111111_1011000111, \
	16'b000000_0011100010, \
	16'b000000_0011001111, \
	16'b111111_1010110110, \
	16'b111111_1111110000, \
	16'b000000_0001110111, \
	16'b000000_0010110110, \
	16'b111111_1101101110, \
	16'b111111_1011011111, \
	16'b111111_1111010011, \
	16'b111111_1101101000, \
	16'b111111_1111000000, \
	16'b111111_1110111110, \
	16'b111111_1110011000, \
	16'b000000_0001101100, \
	16'b000000_0000001111, \
	16'b111111_1111001110, \
	16'b111111_1111101110, \
	16'b000000_0000010100, \
	16'b000000_0000001110, \
	16'b111111_1110011000, \
	16'b111111_1110110100, \
	16'b000000_0001110010, \
	16'b111111_1110101011, \
	16'b111111_1110111101, \
	16'b000000_0001011110, \
	16'b000000_0000100111, \
	16'b111111_1100111000, \
	16'b000000_0001000111, \
	16'b000000_0001001110, \
	16'b000000_0010000100, \
	16'b111111_1111111110, \
	16'b111111_1101010110, \
	16'b000000_0001000000, \
	16'b000000_0001100110, \
	16'b111111_1011000011, \
	16'b111111_1111011010, \
	16'b111111_1111100011, \
	16'b000000_0100011001, \
	16'b111111_1110111001, \
	16'b111111_0110100110, \
	16'b000000_0010010101, \
	16'b000000_0100000111, \
	16'b111111_1001111101, \
	16'b111111_1101110100, \
	16'b000000_0000001110, \
	16'b000000_0100000110, \
	16'b111111_1110010000, \
	16'b111111_1001100011, \
	16'b000000_0001101011, \
	16'b000000_0011001011, \
	16'b111111_1010010101, \
	16'b111111_1110011101, \
	16'b000000_0000111100, \
	16'b000000_0001000111, \
	16'b111111_1111001011, \
	16'b111111_1011010011, \
	16'b000000_0010001110, \
	16'b111111_1111111100, \
	16'b111111_1110001101, \
	16'b111111_1110110001, \
	16'b000000_0000000000, \
	16'b000000_0010000110, \
	16'b111111_1110011110, \
	16'b111111_1101101110, \
	16'b000000_0010001101, \
	16'b111111_1111110001, \
	16'b111111_1111110000, \
	16'b000000_0000001001, \
	16'b111111_1111000111, \
	16'b000000_0010010110, \
	16'b111111_1110000011, \
	16'b000000_0001111000, \
	16'b000000_0010011010, \
	16'b000000_0010000100, \
	16'b000000_0000010001, \
	16'b111111_1110101000, \
	16'b111111_1110010000, \
	16'b000000_0010101010, \
	16'b000000_0000111110, \
	16'b111111_1101100101, \
	16'b000000_0000101110, \
	16'b000000_0001110011, \
	16'b111111_1111110000, \
	16'b000000_0010000001, \
	16'b000000_0000100000, \
	16'b000000_0100101101, \
	16'b111111_1101101001, \
	16'b111111_1001000001, \
	16'b000000_0011100001, \
	16'b000000_0000111010, \
	16'b111111_1101110011, \
	16'b111111_1100100100, \
	16'b000000_0000101010, \
	16'b000000_0100011001, \
	16'b111111_1101100110, \
	16'b111111_1000110100, \
	16'b000000_0010101100, \
	16'b000000_0011011010, \
	16'b111111_1011001111, \
	16'b111111_1110011101, \
	16'b000000_0001001101, \
	16'b000000_0001101000, \
	16'b111111_1111000101, \
	16'b111111_1011001010, \
	16'b000000_0001010000, \
	16'b000000_0000001100, \
	16'b111111_1101101110, \
	16'b111111_1111110110, \
	16'b111111_1110001011, \
	16'b000000_0010011101, \
	16'b111111_1111111100, \
	16'b111111_1111001110, \
	16'b000000_0000101011, \
	16'b111111_1111011100, \
	16'b000000_0000001010, \
	16'b000000_0000100010, \
	16'b000000_0000000111, \
	16'b000000_0001111001, \
	16'b000000_0000000111, \
	16'b000000_0000101011, \
	16'b111111_1111011111, \
	16'b000000_0010011000, \
	16'b111111_1101100110, \
	16'b000000_0001101010, \
	16'b000000_0001101011, \
	16'b000000_0010000000, \
	16'b111111_1111101010, \
	16'b000000_0001100111, \
	16'b000000_0001001010, \
	16'b000000_0010111000, \
	16'b000000_0000000110, \
	16'b111111_1110100100, \
	16'b000000_0000000111, \
	16'b000000_0011111110, \
	16'b111111_1111011000, \
	16'b000000_0001000110, \
	16'b000000_0000111001, \
	16'b000000_0001000101, \
	16'b111111_1101110111, \
	16'b111111_1101110100, \
	16'b000000_0010000001, \
	16'b000000_0011010010, \
	16'b111111_1110110000, \
	16'b000000_0000011101, \
	16'b000000_0010011100, \
	16'b111111_1111100010, \
	16'b111111_1101110110, \
	16'b000000_0000010010, \
	16'b000000_0000000000, \
	16'b000000_0010010110, \
	16'b111111_1110110111, \
	16'b000000_0001100000, \
	16'b000000_0000001100, \
	16'b000000_0001001011, \
	16'b111111_1110100011, \
	16'b111111_1100001000, \
	16'b111111_1101111111, \
	16'b000000_0011001011, \
	16'b000000_0000111001, \
	16'b111111_1111100111, \
	16'b000000_0010110101, \
	16'b000000_0000111000, \
	16'b111111_1110111100, \
	16'b111111_1110101000, \
	16'b000000_0001000111, \
	16'b000000_0000001111, \
	16'b000000_0010000011, \
	16'b111111_1110100110, \
	16'b111111_1110100010, \
	16'b111111_1110011000, \
	16'b000000_0000111110, \
	16'b111111_1110111000, \
	16'b111111_1110111110, \
	16'b111111_1111011101, \
	16'b000000_0000001000, \
	16'b000000_0001000011, \
	16'b111111_1101111100, \
	16'b111111_1100101101, \
	16'b000000_0001001111, \
	16'b111111_1111111111, \
	16'b111111_1110100111, \
	16'b111111_1111001010, \
	16'b111111_1111110110, \
	16'b000000_0001011101, \
	16'b000000_0000111010, \
	16'b111111_1101011111, \
	16'b000000_0010110011, \
	16'b111111_1111110001, \
	16'b111111_1110100110, \
	16'b111111_1111100110, \
	16'b111111_1110111000, \
	16'b000000_0001010001, \
	16'b111111_1110100100, \
	16'b000000_0001010011, \
	16'b000000_0011000111, \
	16'b000000_0001011000, \
	16'b111111_1110000100, \
	16'b111111_1111101010, \
	16'b000000_0001001101, \
	16'b000000_0000000000, \
	16'b111111_1110101100, \
	16'b111111_1111000010, \
	16'b000000_0000101001, \
	16'b000000_0010001100, \
	16'b000000_0001011000, \
	16'b111111_1110101010, \
	16'b111111_1111000011, \
	16'b000000_0000011000, \
	16'b000000_0000000100, \
	16'b000000_0001010011, \
	16'b111111_1111110000, \
	16'b000000_0001100110, \
	16'b000000_0001011101, \
	16'b111111_1110001111, \
	16'b000000_0010101101, \
	16'b000000_0001011100, \
	16'b111111_1110110101, \
	16'b000000_0001100011, \
	16'b111111_1101010011, \
	16'b000000_0000111100, \
	16'b000000_0010010000, \
	16'b111111_1111110101, \
	16'b000000_0001010001, \
	16'b000000_0001101101, \
	16'b111111_1110001001, \
	16'b111111_1101100100, \
	16'b111111_1110011011, \
	16'b000000_0000010000, \
	16'b111111_1111101011, \
	16'b000000_0001000101, \
	16'b111111_1111010110, \
	16'b000000_0000000000, \
	16'b111111_1110001111, \
	16'b111111_1110111110, \
	16'b000000_0100101010, \
	16'b111111_1111001100, \
	16'b111111_1111011101, \
	16'b111111_1110011110, \
	16'b111111_1111110101, \
	16'b111111_1111100100, \
	16'b111111_1111001011, \
	16'b000000_0011011111, \
	16'b000000_0001110100, \
	16'b000000_0010000100, \
	16'b000000_0010000000, \
	16'b111111_1100010111, \
	16'b000000_0010100010, \
	16'b000000_0001110100, \
	16'b111111_1101111100, \
	16'b000000_0100001000, \
	16'b000000_0001011100, \
	16'b000000_0011100100, \
	16'b000000_0001001010, \
	16'b111111_1101110100, \
	16'b000000_0001100011, \
	16'b000000_0000101111, \
	16'b000000_0001011010, \
	16'b000000_0000101010, \
	16'b000000_0001101111, \
	16'b000000_0011110101, \
	16'b000000_0011000111, \
	16'b111111_1110000001, \
	16'b000000_0101100101, \
	16'b111111_1111100001, \
	16'b111111_1111000001, \
	16'b000000_0000001100, \
	16'b000000_0000001001, \
	16'b000000_0011101101, \
	16'b000000_0011010000, \
	16'b000000_0001100000, \
	16'b000000_0001101001, \
	16'b000000_0010101010, \
	16'b000000_0000000100, \
	16'b000000_0010101011, \
	16'b111111_1101011000, \
	16'b000000_0000110000, \
	16'b000000_0001011001, \
	16'b000000_0001110010, \
	16'b111111_1111100110, \
	16'b111111_1110111101, \
	16'b111111_1101101010, \
	16'b000000_0011110110, \
	16'b000000_0000010011, \
	16'b111111_1110100110, \
	16'b111111_1101111000, \
	16'b111111_1101101001, \
	16'b111111_1110001011, \
	16'b111111_1100001110, \
	16'b000000_0010110010, \
	16'b000000_0000101001, \
	16'b111111_1111111101, \
	16'b000000_0000110111, \
	16'b000000_0011010010, \
	16'b111111_1011000101, \
	16'b000000_0001001010, \
	16'b111111_1111011000, \
	16'b000000_0001011011, \
	16'b000000_0100100100, \
	16'b111111_1101101011, \
	16'b000000_0011001100, \
	16'b000000_0101010000, \
	16'b111111_1110011011, \
	16'b000000_0000110110, \
	16'b111111_1011000111, \
	16'b111111_1111110011, \
	16'b000000_0000000000, \
	16'b111111_1110000101, \
	16'b000000_0001011001, \
	16'b000000_0010010010, \
	16'b111111_1101011111, \
	16'b000000_0010100001, \
	16'b111111_1110110110, \
	16'b111111_1111110111, \
	16'b111111_1111011010, \
	16'b111111_1111100000, \
	16'b000000_0101100001, \
	16'b000000_0100110001, \
	16'b111111_1101000010, \
	16'b000000_0010001100, \
	16'b111111_1111010111, \
	16'b000000_0001001010, \
	16'b000000_0010000110, \
	16'b000000_0001111000, \
	16'b000000_0000101011, \
	16'b000000_0010000110, \
	16'b111111_1110101101, \
	16'b111111_1110000101, \
	16'b111111_1111011010, \
	16'b000000_0000011000, \
	16'b000000_0100110010, \
	16'b111111_1110011000, \
	16'b000000_0001101011, \
	16'b111111_1111110000, \
	16'b000000_0000100000, \
	16'b111111_1111100001, \
	16'b000000_0001001001, \
	16'b000000_0010110111, \
	16'b000000_0010001111, \
	16'b111111_1101001110, \
	16'b111111_1111111111, \
	16'b000000_0011110010, \
	16'b111111_1111011110, \
	16'b000000_0011110001, \
	16'b111111_1100101110, \
	16'b000000_0001111001, \
	16'b111111_1110110111, \
	16'b111111_1111110001, \
	16'b000000_0011000100, \
	16'b000000_0110010010, \
	16'b111111_1110101000, \
	16'b000000_0001000100, \
	16'b111111_1111111111, \
	16'b000000_0001111011, \
	16'b111111_1111110101, \
	16'b000000_0001001000, \
	16'b000000_0011001101, \
	16'b000000_0001100001, \
	16'b111111_1110111100, \
	16'b000000_0001110011, \
	16'b000000_0001011000, \
	16'b000000_0000000101, \
	16'b111111_1101110101, \
	16'b000000_0010111100, \
	16'b111111_1111100100, \
	16'b000000_0011101111, \
	16'b111111_1101110000, \
	16'b000000_0001100110, \
	16'b111111_1111101011, \
	16'b111111_1110101111, \
	16'b111111_1111001000, \
	16'b000000_0000100010, \
	16'b000000_0100100011, \
	16'b000000_0001101101, \
	16'b111111_1110100001, \
	16'b111111_1111101010, \
	16'b000000_0000111100, \
	16'b000000_0000111000, \
	16'b000000_1000100001, \
	16'b000000_0001001000, \
	16'b000000_0001110110, \
	16'b000000_0000011100, \
	16'b000000_0001010100, \
	16'b000000_0000010101, \
	16'b000000_0001110011, \
	16'b111111_1111111001, \
	16'b000000_0000110011, \
	16'b111111_1110111100, \
	16'b111111_1111100100, \
	16'b000000_0000000101, \
	16'b000000_0000001000, \
	16'b000000_0010010111, \
	16'b111111_1110101001, \
	16'b000000_0000011000, \
	16'b111111_1100101111, \
	16'b111111_1111100010, \
	16'b000000_0010001011, \
	16'b000000_0010101111, \
	16'b000000_0000000111, \
	16'b000000_0010111000, \
	16'b000000_0000001101, \
	16'b000000_0001010100, \
	16'b111111_1110110000, \
	16'b000000_0000110010, \
	16'b000000_0001110001, \
	16'b111111_1110111010, \
	16'b111111_1110101011, \
	16'b000000_0000010110, \
	16'b111111_1110010100, \
	16'b111111_1110111111, \
	16'b000000_0000100001, \
	16'b000000_0001010110, \
	16'b000000_0001001110, \
	16'b000000_0000101000, \
	16'b111111_1110011111, \
	16'b000000_0000110010, \
	16'b111111_1111110000, \
	16'b111111_1101110100, \
	16'b111111_1111110000, \
	16'b000000_0001110111, \
	16'b000000_0010110010, \
	16'b111111_1110000111, \
	16'b111111_1111010111, \
	16'b111111_1111001110, \
	16'b000000_0000011000, \
	16'b111111_1111000111, \
	16'b111111_1101101010, \
	16'b111111_1111000111, \
	16'b000000_0010100010, \
	16'b000000_0000100110, \
	16'b111111_1110100010, \
	16'b000000_0001101000, \
	16'b111111_1110001011, \
	16'b111111_1111001100, \
	16'b111111_1110100000, \
	16'b111111_1111101001, \
	16'b000000_0001111111, \
	16'b000000_0001010100, \
	16'b000000_0000010110, \
	16'b000000_0010101010, \
	16'b111111_1111000100, \
	16'b000000_0000101010, \
	16'b111111_1111011101, \
	16'b000000_0000111101, \
	16'b000000_0010011010, \
	16'b000000_0000111111, \
	16'b111111_1111100110, \
	16'b000000_0001000011, \
	16'b111111_1110100110, \
	16'b000000_0000001111, \
	16'b000000_0000011001, \
	16'b111111_1111100011, \
	16'b000000_0010011001, \
	16'b000000_0000010011\
};

`define maxpool_biases_PDMHN parameter bit [15:0] maxpool_biases_PDMHN [9:0] = '{ \
	16'b111111_1110101110, \
	16'b111111_1001010001, \
	16'b000000_0011010010, \
	16'b111111_1111100000, \
	16'b111111_1111100010, \
	16'b000000_0000001111, \
	16'b111111_1100110011, \
	16'b000000_0001001011, \
	16'b000000_1001010101, \
	16'b111111_1110001100\
};

module Maxpool_FC_YJWNR(
	input    clk,
	input    reset,
	input    valid,
	output reg   done,
	output reg   ready,
	output reg  [10:0] inp_addr,
	input   [15:0] inp_data,
	output reg  [3:0] out_addr,
	output reg  [15:0] out_data,
	output reg   out_we
);
	`maxpool_weights_JWCVA
	`maxpool_biases_PDMHN

	reg  [11:0] weights_ra;
	wire  [15:0] weights_rd;
	reg  [3:0] biases_ra;
	wire  [15:0] biases_rd;
	reg signed [15:0] window [31:0];
	reg signed [15:0] mp_out [287:0];
	reg  [10:0] curr_y;
	reg  [8:0] out_y;
	reg  [10:0] curr_x;
	reg  [8:0] out_x;
	reg  [10:0] jj;
	reg  [10:0] ii;
	reg  [10:0] kk;
	reg  [4:0] ww;
	reg  [3:0] wc;
	reg  [4:0] wr;
	wire signed [15:0] max_out;
	wire signed [15:0] max_logic_VDSRS;
	wire signed [15:0] max_logic_CCYVZ;
	wire signed [15:0] max_logic_HIGIY;
	wire signed [15:0] max_logic_JPOTC;
	wire signed [15:0] max_logic_SRNNQ;
	wire signed [15:0] max_logic_HGNVV;
	wire signed [15:0] max_logic_NQMVI;
	wire signed [15:0] max_logic_BRCGE;
	wire signed [15:0] max_logic_WASXX;
	wire signed [15:0] max_logic_UYMTD;
	wire signed [15:0] max_logic_URZFO;
	wire signed [15:0] max_logic_QBPPZ;
	wire signed [15:0] max_logic_GLWCV;
	wire signed [15:0] max_logic_TKYYU;
	wire signed [15:0] max_logic_AVFGO;
	wire signed [15:0] max_logic_CSGPI;
	wire signed [15:0] max_logic_ZZGYI;
	wire signed [15:0] max_logic_LKYAV;
	wire signed [15:0] max_logic_BTFOH;
	wire signed [15:0] max_logic_DOROX;
	wire signed [15:0] max_logic_ZQGMQ;
	wire signed [15:0] max_logic_MOZBT;
	wire signed [15:0] max_logic_ILWCY;
	wire signed [15:0] max_logic_BEULH;
	reg signed [15:0] dot_product;
	wire signed [15:0] prod;
	reg  [3:0] state;


	// tie the weight data to the weight address
	assign weights_rd = maxpool_weights_JWCVA[weights_ra];

	// tie the bias data to the bias address
	assign biases_rd = maxpool_biases_PDMHN[biases_ra];

	// instantiate the state machine
	always @ (posedge clk) begin
		if (reset) begin
			// clear done flag and go to starting state
			done <= 1'd0;
			inp_addr <= 11'd0;
			weights_ra <= 12'd0;
			biases_ra <= 4'd0;
			out_addr <= 4'd0;
			out_we <= 1'd0;
			curr_y <= 11'd0;
			out_y <= 9'd0;
			curr_x <= 11'd0;
			out_x <= 9'd0;
			dot_product <= 16'd0;
			state <= 4'd0;
		end
		else begin
			case (state)
				// _StWaitValid
				4'd0: begin
						if (valid) begin
							state <= 4'd1;
						end
					end
				// _StResetWindow
				4'd1: begin
						jj <= 11'd0;
						ii <= 11'd0;
						kk <= 11'd0;
						ww <= 5'd0;
						state <= 4'd2;
					end
				// _StSetInpAddr
				4'd2: begin
						inp_addr <= (curr_y + jj) * 11'd12 * 11'd8 + (curr_x + ii) * 11'd8 + kk;
						state <= 4'd3;
					end
				// _StWindowBuffer
				4'd3: begin
						state <= 4'd4;
					end
				// _StSetWindow
				4'd4: begin
						window[ww] <= inp_data;
						if (ww == 5'd31) begin
							state <= 4'd5;
						end
						else begin
							ww <= ww + 5'd1;
							if (kk == 11'd7) begin
								kk <= 11'd0;
								if (ii == 11'd1) begin
									ii <= 11'd0;
									jj <= jj + 11'd1;
								end
								else begin
									ii <= ii + 11'd1;
								end
							end
							else begin
								kk <= kk + 11'd1;
							end
							state <= 4'd2;
						end
					end
				// _StFindMax
				4'd5: begin
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd0] <= max_logic_HIGIY;
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd1] <= max_logic_HGNVV;
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd2] <= max_logic_WASXX;
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd3] <= max_logic_QBPPZ;
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd4] <= max_logic_AVFGO;
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd5] <= max_logic_LKYAV;
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd6] <= max_logic_ZQGMQ;
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd7] <= max_logic_BEULH;
						state <= 4'd6;
					end
				// _StIncMaxpool
				4'd6: begin
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd0] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd0];
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd1] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd1];
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd2] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd2];
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd3] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd3];
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd4] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd4];
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd5] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd5];
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd6] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd6];
						mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd7] <= mp_out[out_y * 9'd6 * 9'd8 + out_x * 9'd8 + 9'd7];
						if (curr_x > 11'd8) begin
							curr_x <= 11'd0;
							out_x <= 9'd0;
							if (curr_y > 11'd8) begin
								state <= 4'd7;
							end
							else begin
								curr_y <= curr_y + 11'd2;
								out_y <= out_y + 9'd1;
								state <= 4'd1;
							end
						end
						else begin
							curr_x <= curr_x + 11'd2;
							out_x <= out_x + 9'd1;
							state <= 4'd1;
						end
					end
				// _StWaitDotProduct
				4'd7: begin
						dot_product <= dot_product + prod;
						

						if (out_x == 9'd287) begin
							weights_ra <= weights_ra + 12'd1;
							out_we <= 1'd1;
							out_data <= dot_product + prod + maxpool_biases_PDMHN[out_addr];
							state <= 4'd8;
						end
						else begin
							out_x <= out_x + 9'd1;
							weights_ra <= weights_ra + 12'd1;
						end
					end
				// _StWriteData
				4'd8: begin
						out_we <= 1'd0;
						out_x <= 9'd0;
						dot_product <= 16'd0;
						if (out_addr == 9) begin
							state <= 4'd9;
						end
						else begin
							out_addr <= out_addr + 4'd1;
							state <= 4'd7;
						end
					end
				// V_StDone
				4'd9: begin
						// idle until reset
						done <= 1'd1;
						state <= 4'd9;
					end
			endcase
		end
	end
	// instantiate the signed maximum modules
	SignedMax_RRWYK SignedMax_RRWYK_VKNLU(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[0]), 
		.input_SWLTH(window[8]), 
		.output_MHDGF(max_logic_VDSRS)
	);

	SignedMax_RRWYK SignedMax_RRWYK_EIKYH(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[16]), 
		.input_SWLTH(window[24]), 
		.output_MHDGF(max_logic_CCYVZ)
	);

	SignedMax_RRWYK SignedMax_RRWYK_EAUUN(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_VDSRS), 
		.input_SWLTH(max_logic_CCYVZ), 
		.output_MHDGF(max_logic_HIGIY)
	);

	SignedMax_RRWYK SignedMax_RRWYK_WVCSV(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[1]), 
		.input_SWLTH(window[9]), 
		.output_MHDGF(max_logic_JPOTC)
	);

	SignedMax_RRWYK SignedMax_RRWYK_ZNEXX(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[17]), 
		.input_SWLTH(window[25]), 
		.output_MHDGF(max_logic_SRNNQ)
	);

	SignedMax_RRWYK SignedMax_RRWYK_VEZHK(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_JPOTC), 
		.input_SWLTH(max_logic_SRNNQ), 
		.output_MHDGF(max_logic_HGNVV)
	);

	SignedMax_RRWYK SignedMax_RRWYK_CPVXI(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[2]), 
		.input_SWLTH(window[10]), 
		.output_MHDGF(max_logic_NQMVI)
	);

	SignedMax_RRWYK SignedMax_RRWYK_MELAM(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[18]), 
		.input_SWLTH(window[26]), 
		.output_MHDGF(max_logic_BRCGE)
	);

	SignedMax_RRWYK SignedMax_RRWYK_BVJHX(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_NQMVI), 
		.input_SWLTH(max_logic_BRCGE), 
		.output_MHDGF(max_logic_WASXX)
	);

	SignedMax_RRWYK SignedMax_RRWYK_DYDPU(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[3]), 
		.input_SWLTH(window[11]), 
		.output_MHDGF(max_logic_UYMTD)
	);

	SignedMax_RRWYK SignedMax_RRWYK_CXYIP(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[19]), 
		.input_SWLTH(window[27]), 
		.output_MHDGF(max_logic_URZFO)
	);

	SignedMax_RRWYK SignedMax_RRWYK_OXCQM(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_UYMTD), 
		.input_SWLTH(max_logic_URZFO), 
		.output_MHDGF(max_logic_QBPPZ)
	);

	SignedMax_RRWYK SignedMax_RRWYK_SZQLP(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[4]), 
		.input_SWLTH(window[12]), 
		.output_MHDGF(max_logic_GLWCV)
	);

	SignedMax_RRWYK SignedMax_RRWYK_GFGZG(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[20]), 
		.input_SWLTH(window[28]), 
		.output_MHDGF(max_logic_TKYYU)
	);

	SignedMax_RRWYK SignedMax_RRWYK_TGMBV(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_GLWCV), 
		.input_SWLTH(max_logic_TKYYU), 
		.output_MHDGF(max_logic_AVFGO)
	);

	SignedMax_RRWYK SignedMax_RRWYK_ZVMBI(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[5]), 
		.input_SWLTH(window[13]), 
		.output_MHDGF(max_logic_CSGPI)
	);

	SignedMax_RRWYK SignedMax_RRWYK_GACAF(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[21]), 
		.input_SWLTH(window[29]), 
		.output_MHDGF(max_logic_ZZGYI)
	);

	SignedMax_RRWYK SignedMax_RRWYK_ZVDAL(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_CSGPI), 
		.input_SWLTH(max_logic_ZZGYI), 
		.output_MHDGF(max_logic_LKYAV)
	);

	SignedMax_RRWYK SignedMax_RRWYK_QLSIY(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[6]), 
		.input_SWLTH(window[14]), 
		.output_MHDGF(max_logic_BTFOH)
	);

	SignedMax_RRWYK SignedMax_RRWYK_FGHDZ(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[22]), 
		.input_SWLTH(window[30]), 
		.output_MHDGF(max_logic_DOROX)
	);

	SignedMax_RRWYK SignedMax_RRWYK_DCJXE(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_BTFOH), 
		.input_SWLTH(max_logic_DOROX), 
		.output_MHDGF(max_logic_ZQGMQ)
	);

	SignedMax_RRWYK SignedMax_RRWYK_OANZE(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[7]), 
		.input_SWLTH(window[15]), 
		.output_MHDGF(max_logic_MOZBT)
	);

	SignedMax_RRWYK SignedMax_RRWYK_YHALR(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(window[23]), 
		.input_SWLTH(window[31]), 
		.output_MHDGF(max_logic_ILWCY)
	);

	SignedMax_RRWYK SignedMax_RRWYK_XCBQQ(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_HKTGS(max_logic_MOZBT), 
		.input_SWLTH(max_logic_ILWCY), 
		.output_MHDGF(max_logic_BEULH)
	);


	// instantiate the multiplier
	SignedMult_MRMTA SignedMult_MRMTA_OPXHL(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_TUOCE(mp_out[out_x]), 
		.input_IXGYP(weights_rd), 
		.output_XWLZX(prod)
	);


endmodule



module SignedMax_RRWYK(
	input    clk,
	input    reset,
	input    valid,
	output    done,
	output reg   ready,
	input  signed [15:0] input_HKTGS,
	input  signed [15:0] input_SWLTH,
	output  signed [15:0] output_MHDGF
);


	// tie `done` to `HIGH`
	assign done = 1'd1;

	// use ternary to determine the max
	assign output_MHDGF = (input_HKTGS > input_SWLTH) ? 
		input_HKTGS : 
		input_SWLTH;

endmodule



module SignedMult_MRMTA(
	input    clk,
	input    reset,
	input    valid,
	output    done,
	output reg   ready,
	input  signed [15:0] input_TUOCE,
	input  signed [15:0] input_IXGYP,
	output  signed [15:0] output_XWLZX
);

	wire signed [31:0] mult_out;

	// tie `done` to `HIGH`
	assign done = 1'd1;

	// intermediate full bit length mult
	assign mult_out = input_TUOCE * input_IXGYP;

	// select bits for `N.M` fixed point
	assign output_XWLZX = {mult_out[31], mult_out[24:10]};

endmodule



`endif