// synthesis VERILOG_INPUT_VERSION SYSTEMVERILOG_2005
`ifndef __LAYER3_SV__
`define __LAYER3_SV__



`define conv2dsum1d_weights_KLAOE parameter bit [15:0] conv2dsum1d_weights_KLAOE [255:0] = '{ \
	16'b111111_1100001010, \
	16'b000000_0111100010, \
	16'b000000_0010110011, \
	16'b111111_1011111010, \
	16'b000000_0101100001, \
	16'b000000_1000101100, \
	16'b000000_0111101000, \
	16'b000000_0001011101, \
	16'b000000_0001110011, \
	16'b000000_0011101100, \
	16'b111111_1111111110, \
	16'b000000_0011110010, \
	16'b111111_1111010100, \
	16'b111111_1110111001, \
	16'b000000_0010001011, \
	16'b000000_0101110011, \
	16'b000000_0010110000, \
	16'b111110_1011100110, \
	16'b111111_1011101000, \
	16'b111111_1100101001, \
	16'b111111_0000001110, \
	16'b111111_1000100111, \
	16'b111111_0111010001, \
	16'b111111_1010100000, \
	16'b111111_1011110011, \
	16'b111111_0111101100, \
	16'b000000_0010111101, \
	16'b111111_1100000111, \
	16'b111111_1011100000, \
	16'b000000_0000010000, \
	16'b111111_1100000111, \
	16'b111111_1111110010, \
	16'b111111_1111011001, \
	16'b111111_0010110010, \
	16'b111111_1010111100, \
	16'b111111_1010010100, \
	16'b111111_1010011010, \
	16'b000000_0010001011, \
	16'b111111_1100010000, \
	16'b111111_1110010101, \
	16'b000000_0011010101, \
	16'b000000_1101101000, \
	16'b000000_0010000100, \
	16'b000000_0011100100, \
	16'b000000_0111001111, \
	16'b000000_0000110000, \
	16'b000000_1001001111, \
	16'b111111_1010100100, \
	16'b000000_0100011010, \
	16'b000000_1101011101, \
	16'b000000_0100011101, \
	16'b000000_0001100100, \
	16'b000000_1010110110, \
	16'b111111_1110000001, \
	16'b000000_0010011111, \
	16'b000000_1000111101, \
	16'b000000_0001101000, \
	16'b111111_0110100001, \
	16'b111111_1110101110, \
	16'b111111_1100100000, \
	16'b111111_0011110001, \
	16'b111111_1000110110, \
	16'b111111_1100010010, \
	16'b111111_1000001011, \
	16'b000000_0011101101, \
	16'b111111_0011100110, \
	16'b000000_0011000101, \
	16'b111111_1010000001, \
	16'b111111_1010110010, \
	16'b000000_0011000011, \
	16'b111111_1001110110, \
	16'b111111_0110101101, \
	16'b000000_0011110100, \
	16'b000000_1011110100, \
	16'b000000_0000010011, \
	16'b000000_0111111010, \
	16'b000000_1101000101, \
	16'b000000_0000111100, \
	16'b111111_1110101000, \
	16'b000000_1011001010, \
	16'b111111_1111111000, \
	16'b111110_1110000001, \
	16'b000000_0001001111, \
	16'b111111_1011010110, \
	16'b111111_0110010011, \
	16'b111111_1100010100, \
	16'b111111_1010010011, \
	16'b111111_1000011010, \
	16'b111111_1011101011, \
	16'b111111_1111011010, \
	16'b000000_0101000000, \
	16'b111111_1111001101, \
	16'b000000_0110000100, \
	16'b000000_0101110000, \
	16'b000000_0100001011, \
	16'b000000_0101001000, \
	16'b111111_1111111000, \
	16'b111111_0110001011, \
	16'b111111_1011101111, \
	16'b111111_1111000111, \
	16'b111111_1110110011, \
	16'b111111_1101001101, \
	16'b111111_1100011010, \
	16'b111111_1010000000, \
	16'b000000_0100011010, \
	16'b000001_0010011011, \
	16'b111111_1101001001, \
	16'b000000_0100100111, \
	16'b000000_1101101111, \
	16'b000000_0001001101, \
	16'b000000_1000110011, \
	16'b000000_0000011101, \
	16'b000000_0011010100, \
	16'b111111_0100110110, \
	16'b000000_0000110010, \
	16'b111111_1011100011, \
	16'b000000_0000000011, \
	16'b111111_1100000011, \
	16'b111111_0110101110, \
	16'b000000_0000001110, \
	16'b000000_0100110101, \
	16'b000000_1110101011, \
	16'b000000_0111101110, \
	16'b000000_0010001011, \
	16'b000000_1011000110, \
	16'b000000_0110101000, \
	16'b000000_0101001110, \
	16'b000000_1001100010, \
	16'b000000_0010111100, \
	16'b111111_0001100110, \
	16'b111111_1010010111, \
	16'b111111_1100010111, \
	16'b111111_0111010010, \
	16'b111111_1101110011, \
	16'b000000_0001001110, \
	16'b111111_0011110001, \
	16'b111111_1100001110, \
	16'b000000_0111000011, \
	16'b000000_0011001100, \
	16'b000000_0010111111, \
	16'b000000_0110000011, \
	16'b111111_1010001110, \
	16'b111111_1011010001, \
	16'b000000_1001101110, \
	16'b000000_0110101010, \
	16'b000000_1100010000, \
	16'b111111_1001101110, \
	16'b111111_1100101101, \
	16'b000000_0111010001, \
	16'b000000_0001000001, \
	16'b000000_0100001010, \
	16'b000000_1110100101, \
	16'b000000_0001100010, \
	16'b111111_1100010110, \
	16'b111111_1101000000, \
	16'b111111_1110101101, \
	16'b111111_1010110101, \
	16'b000000_0001100101, \
	16'b111111_1100110000, \
	16'b111111_1010011000, \
	16'b111111_1111111001, \
	16'b000000_0100000001, \
	16'b000000_0100100111, \
	16'b000000_0011001011, \
	16'b000000_1101000111, \
	16'b000000_0010111100, \
	16'b000000_0110100011, \
	16'b000000_1111000100, \
	16'b111111_1110110010, \
	16'b111111_0010001010, \
	16'b111111_1011001111, \
	16'b000000_0010110101, \
	16'b111111_0110000111, \
	16'b111111_1010001111, \
	16'b111111_0110110001, \
	16'b111111_0011010101, \
	16'b000000_0000111000, \
	16'b000000_0011000100, \
	16'b000000_0000110000, \
	16'b000000_0011001011, \
	16'b000000_0011111011, \
	16'b111111_1001111101, \
	16'b111111_1101101111, \
	16'b000000_0101111011, \
	16'b111111_1111001101, \
	16'b111111_1001101001, \
	16'b000000_0011011010, \
	16'b111111_1011101010, \
	16'b111111_0110111110, \
	16'b111111_0110100011, \
	16'b111111_1100101100, \
	16'b111111_1110110110, \
	16'b111111_1011000010, \
	16'b111111_1001001101, \
	16'b111111_1011111110, \
	16'b111111_1101000001, \
	16'b111111_1100000010, \
	16'b000000_0100101100, \
	16'b000000_0011011001, \
	16'b000000_0100111011, \
	16'b111111_1011110101, \
	16'b111111_1011100001, \
	16'b111111_1110001001, \
	16'b111111_1101100110, \
	16'b000000_0000110001, \
	16'b111111_1011010011, \
	16'b111111_1001101110, \
	16'b000000_0101110001, \
	16'b000000_0000110101, \
	16'b000000_1100110000, \
	16'b111111_1100000111, \
	16'b000000_0101001010, \
	16'b000000_0100111101, \
	16'b000000_0001110100, \
	16'b000000_1011101100, \
	16'b000000_1011111010, \
	16'b000000_0011010111, \
	16'b111111_1100101010, \
	16'b000000_0000010111, \
	16'b111111_1100110011, \
	16'b000000_0101001111, \
	16'b000000_0011100010, \
	16'b000000_0010011000, \
	16'b000000_0000001100, \
	16'b000000_0011100011, \
	16'b111111_1000011110, \
	16'b111111_1011100010, \
	16'b111111_1111011111, \
	16'b111111_0110010000, \
	16'b000000_0010110111, \
	16'b111111_1100100101, \
	16'b111111_0111010100, \
	16'b111111_1111010100, \
	16'b111110_1101111100, \
	16'b111111_1111010111, \
	16'b111111_0111100011, \
	16'b111111_0101101011, \
	16'b000000_0001101001, \
	16'b111111_1000100011, \
	16'b111111_0001010100, \
	16'b000000_0100111110, \
	16'b000000_1100000011, \
	16'b000000_0010010001, \
	16'b111111_1110111011, \
	16'b000000_1001101001, \
	16'b111111_1010101010, \
	16'b111111_1010000110, \
	16'b000000_1010110001, \
	16'b000000_0011001010, \
	16'b000000_1010110110, \
	16'b000000_0110001111, \
	16'b000000_0110111110, \
	16'b000000_0110001101, \
	16'b000000_0000111110, \
	16'b111111_1111010011, \
	16'b000000_0101001000\
};

`define conv2dsum1d_biases_USXDE parameter bit [15:0] conv2dsum1d_biases_USXDE [7:0] = '{ \
	16'b000000_1011001100, \
	16'b111111_1000010100, \
	16'b000000_0101010010, \
	16'b000000_0010011100, \
	16'b000000_0011010101, \
	16'b000000_0000010000, \
	16'b111111_0100110000, \
	16'b111111_1100110011\
};

module Conv2DSum1D_LXJTZ(
	input    clk,
	input    reset,
	input    valid,
	output reg   done,
	output reg   ready,
	output reg  [10:0] inp_addr,
	input  signed [15:0] inp_data,
	output reg  [10:0] out_addr,
	output reg  [15:0] out_data,
	output reg   out_we
);
	`conv2dsum1d_weights_KLAOE
	`conv2dsum1d_biases_USXDE

	reg  [7:0] weights_ra;
	wire  [15:0] weights_rd;
	reg  [2:0] biases_ra;
	wire  [15:0] biases_rd;
	reg  [10:0] ti;
	reg  [10:0] tj;
	reg  [7:0] wc;
	reg  [10:0] cr;
	reg  [13:0] oc;
	reg  [10:0] ii;
	reg  [10:0] jj;
	reg  [10:0] r;
	reg signed [15:0] sub_img [3:0];
	reg signed [15:0] sum_arr [7:0];
	wire signed [15:0] mult_out_0;
	wire signed [15:0] mult_out_1;
	wire signed [15:0] mult_out_2;
	wire signed [15:0] mult_out_3;
	reg  [3:0] state;


	// tie the weight data to the weight address
	assign weights_rd = conv2dsum1d_weights_KLAOE[weights_ra];

	// tie the bias data to the bias address
	assign biases_rd = conv2dsum1d_biases_USXDE[biases_ra];

	// instantiate the state machine
	always @ (posedge clk) begin
		if (reset) begin
			// clear done flag and go to starting state
			done <= 1'd0;
			inp_addr <= 11'd0;
			biases_ra <= 3'd0;
			out_addr <= 11'd0;
			out_we <= 1'd0;
			ti <= 11'd0;
			tj <= 11'd0;
			wc <= 8'd0;
			cr <= 11'd0;
			oc <= 14'd0;
			state <= 4'd0;
		end
		else begin
			case (state)
				// _StWaitValid
				4'd0: begin
						if (valid) begin
							state <= 4'd1;
						end
					end
				// _StResetSumArr
				4'd1: begin
						sum_arr[0] <= 16'd0;
						sum_arr[1] <= 16'd0;
						sum_arr[2] <= 16'd0;
						sum_arr[3] <= 16'd0;
						sum_arr[4] <= 16'd0;
						sum_arr[5] <= 16'd0;
						sum_arr[6] <= 16'd0;
						sum_arr[7] <= 16'd0;
						state <= 4'd2;
					end
				// _StResetSub
				4'd2: begin
						ii <= 11'd0;
						jj <= 11'd0;
						r <= 11'd0;
						state <= 4'd3;
					end
				// _StSetInpAddr
				4'd3: begin
						inp_addr <= (ti + ii) * 11'd13 * 11'd8 + (tj + jj) * 11'd8 + cr;
						state <= 4'd4;
					end
				// _StSubBuffer
				4'd4: begin
						state <= 4'd5;
					end
				// _StSetSub
				4'd5: begin
						sub_img[r] <= inp_data;
						if (r == 11'd3) begin
							wc <= 8'd0;
							state <= 4'd6;
						end
						else begin
							r <= r + 11'd1;
							if (jj == 11'd1) begin
								ii <= ii + 11'd1;
								jj <= 11'd0;
							end
							else begin
								jj <= jj + 11'd1;
							end
							state <= 4'd3;
						end
					end
				// _StComputeConv
				4'd6: begin
						// assign the output of the convolution
						sum_arr[wc] <= sum_arr[wc] + 
		mult_out_0 + 
		mult_out_1 + 
		mult_out_2 + 
		mult_out_3;
						state <= 4'd7;
					end
				// _StIncWeightIndices
				4'd7: begin
						if (wc == 8'd7) begin
							wc <= 8'd0;
							if (oc == 14'd9215) begin
								oc <= 14'd0;
								state <= 4'd8;
							end
							else begin
								oc <= oc + 14'd1;
								state <= 4'd8;
							end
						end
						else begin
							wc <= wc + 8'd1;
							oc <= oc + 14'd1;
							state <= 4'd6;
						end
					end
				// _StIncTargetIndices
				4'd8: begin
						if (cr == 11'd7) begin
							cr <= 11'd0;
							if (tj == 11'd11) begin
								tj <= 11'd0;
								if (ti == 11'd11) begin
									ti <= 11'd0;
								end
								else begin
									ti <= ti + 11'd1;
								end
							end
							else begin
								tj <= tj + 11'd1;
							end
							state <= 4'd9;
						end
						else begin
							cr <= cr + 11'd1;
							state <= 4'd2;
						end
					end
				// _StWriteData
				4'd9: begin
						out_data <= sum_arr[wc] + conv2dsum1d_biases_USXDE[wc];
						if (out_addr == 1152) begin
							state <= 4'd11;
						end
						else begin
							if (wc == 8'd8) begin
								wc <= 8'd0;
								state <= 4'd1;
							end
							else begin
								out_we <= 1'd1;
								state <= 4'd10;
							end
						end
					end
				// _StWriteBuffer
				4'd10: begin
						out_we <= 1'd0;
						out_addr <= out_addr + 11'd1;
						wc <= wc + 8'd1;
						state <= 4'd9;
					end
				// V_StDone
				4'd11: begin
						// idle until reset
						done <= 1'd1;
						state <= 4'd11;
					end
			endcase
		end
	end
	// instantiate the multipliers
	SignedMult_FAIDC SignedMult_FAIDC_JCNFX(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_AEOFK(sub_img[0]), 
		.input_KMKQK(conv2dsum1d_weights_KLAOE[wc * 8'd8 + cr + 8'd0]), 
		.output_OCNPV(mult_out_0)
	);

	SignedMult_FAIDC SignedMult_FAIDC_TXHYV(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_AEOFK(sub_img[1]), 
		.input_KMKQK(conv2dsum1d_weights_KLAOE[wc * 8'd8 + cr + 8'd64]), 
		.output_OCNPV(mult_out_1)
	);

	SignedMult_FAIDC SignedMult_FAIDC_MWWSL(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_AEOFK(sub_img[2]), 
		.input_KMKQK(conv2dsum1d_weights_KLAOE[wc * 8'd8 + cr + 8'd128]), 
		.output_OCNPV(mult_out_2)
	);

	SignedMult_FAIDC SignedMult_FAIDC_JOBVH(
		.clk(), 
		.reset(), 
		.valid(), 
		.done(), 
		.ready(), 
		.input_AEOFK(sub_img[3]), 
		.input_KMKQK(conv2dsum1d_weights_KLAOE[wc * 8'd8 + cr + 8'd192]), 
		.output_OCNPV(mult_out_3)
	);


endmodule



module SignedMult_FAIDC(
	input    clk,
	input    reset,
	input    valid,
	output    done,
	output reg   ready,
	input  signed [15:0] input_AEOFK,
	input  signed [15:0] input_KMKQK,
	output  signed [15:0] output_OCNPV
);

	wire signed [31:0] mult_out;

	// tie `done` to `HIGH`
	assign done = 1'd1;

	// intermediate full bit length mult
	assign mult_out = input_AEOFK * input_KMKQK;

	// select bits for `N.M` fixed point
	assign output_OCNPV = {mult_out[31], mult_out[24:10]};

endmodule



`endif